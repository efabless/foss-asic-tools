magic
tech sky130A
magscale 1 2
timestamp 1374899056
<< checkpaint >>
rect -1139 -1208 2343 3918
<< pwell >>
rect 215 2382 989 2658
rect 121 1612 1083 1874
rect 121 436 1083 698
<< nmos >>
rect 200 1638 230 1848
rect 286 1638 316 1848
rect 372 1638 402 1848
rect 458 1638 488 1848
rect 544 1638 574 1848
rect 630 1638 660 1848
rect 716 1638 746 1848
rect 802 1638 832 1848
rect 888 1638 918 1848
rect 974 1638 1004 1848
rect 200 462 230 672
rect 286 462 316 672
rect 372 462 402 672
rect 458 462 488 672
rect 544 462 574 672
rect 630 462 660 672
rect 716 462 746 672
rect 802 462 832 672
rect 888 462 918 672
rect 974 462 1004 672
<< ndiff >>
rect 147 1824 200 1848
rect 147 1790 155 1824
rect 189 1790 200 1824
rect 147 1756 200 1790
rect 147 1722 155 1756
rect 189 1722 200 1756
rect 147 1688 200 1722
rect 147 1654 155 1688
rect 189 1654 200 1688
rect 147 1638 200 1654
rect 230 1824 286 1848
rect 230 1790 241 1824
rect 275 1790 286 1824
rect 230 1756 286 1790
rect 230 1722 241 1756
rect 275 1722 286 1756
rect 230 1688 286 1722
rect 230 1654 241 1688
rect 275 1654 286 1688
rect 230 1638 286 1654
rect 316 1824 372 1848
rect 316 1790 327 1824
rect 361 1790 372 1824
rect 316 1756 372 1790
rect 316 1722 327 1756
rect 361 1722 372 1756
rect 316 1688 372 1722
rect 316 1654 327 1688
rect 361 1654 372 1688
rect 316 1638 372 1654
rect 402 1824 458 1848
rect 402 1790 413 1824
rect 447 1790 458 1824
rect 402 1756 458 1790
rect 402 1722 413 1756
rect 447 1722 458 1756
rect 402 1688 458 1722
rect 402 1654 413 1688
rect 447 1654 458 1688
rect 402 1638 458 1654
rect 488 1824 544 1848
rect 488 1790 499 1824
rect 533 1790 544 1824
rect 488 1756 544 1790
rect 488 1722 499 1756
rect 533 1722 544 1756
rect 488 1688 544 1722
rect 488 1654 499 1688
rect 533 1654 544 1688
rect 488 1638 544 1654
rect 574 1824 630 1848
rect 574 1790 585 1824
rect 619 1790 630 1824
rect 574 1756 630 1790
rect 574 1722 585 1756
rect 619 1722 630 1756
rect 574 1688 630 1722
rect 574 1654 585 1688
rect 619 1654 630 1688
rect 574 1638 630 1654
rect 660 1824 716 1848
rect 660 1790 671 1824
rect 705 1790 716 1824
rect 660 1756 716 1790
rect 660 1722 671 1756
rect 705 1722 716 1756
rect 660 1688 716 1722
rect 660 1654 671 1688
rect 705 1654 716 1688
rect 660 1638 716 1654
rect 746 1824 802 1848
rect 746 1790 757 1824
rect 791 1790 802 1824
rect 746 1756 802 1790
rect 746 1722 757 1756
rect 791 1722 802 1756
rect 746 1688 802 1722
rect 746 1654 757 1688
rect 791 1654 802 1688
rect 746 1638 802 1654
rect 832 1824 888 1848
rect 832 1790 843 1824
rect 877 1790 888 1824
rect 832 1756 888 1790
rect 832 1722 843 1756
rect 877 1722 888 1756
rect 832 1688 888 1722
rect 832 1654 843 1688
rect 877 1654 888 1688
rect 832 1638 888 1654
rect 918 1824 974 1848
rect 918 1790 929 1824
rect 963 1790 974 1824
rect 918 1756 974 1790
rect 918 1722 929 1756
rect 963 1722 974 1756
rect 918 1688 974 1722
rect 918 1654 929 1688
rect 963 1654 974 1688
rect 918 1638 974 1654
rect 1004 1824 1057 1848
rect 1004 1790 1015 1824
rect 1049 1790 1057 1824
rect 1004 1756 1057 1790
rect 1004 1722 1015 1756
rect 1049 1722 1057 1756
rect 1004 1688 1057 1722
rect 1004 1654 1015 1688
rect 1049 1654 1057 1688
rect 1004 1638 1057 1654
rect 147 648 200 672
rect 147 614 155 648
rect 189 614 200 648
rect 147 580 200 614
rect 147 546 155 580
rect 189 546 200 580
rect 147 512 200 546
rect 147 478 155 512
rect 189 478 200 512
rect 147 462 200 478
rect 230 648 286 672
rect 230 614 241 648
rect 275 614 286 648
rect 230 580 286 614
rect 230 546 241 580
rect 275 546 286 580
rect 230 512 286 546
rect 230 478 241 512
rect 275 478 286 512
rect 230 462 286 478
rect 316 648 372 672
rect 316 614 327 648
rect 361 614 372 648
rect 316 580 372 614
rect 316 546 327 580
rect 361 546 372 580
rect 316 512 372 546
rect 316 478 327 512
rect 361 478 372 512
rect 316 462 372 478
rect 402 648 458 672
rect 402 614 413 648
rect 447 614 458 648
rect 402 580 458 614
rect 402 546 413 580
rect 447 546 458 580
rect 402 512 458 546
rect 402 478 413 512
rect 447 478 458 512
rect 402 462 458 478
rect 488 648 544 672
rect 488 614 499 648
rect 533 614 544 648
rect 488 580 544 614
rect 488 546 499 580
rect 533 546 544 580
rect 488 512 544 546
rect 488 478 499 512
rect 533 478 544 512
rect 488 462 544 478
rect 574 648 630 672
rect 574 614 585 648
rect 619 614 630 648
rect 574 580 630 614
rect 574 546 585 580
rect 619 546 630 580
rect 574 512 630 546
rect 574 478 585 512
rect 619 478 630 512
rect 574 462 630 478
rect 660 648 716 672
rect 660 614 671 648
rect 705 614 716 648
rect 660 580 716 614
rect 660 546 671 580
rect 705 546 716 580
rect 660 512 716 546
rect 660 478 671 512
rect 705 478 716 512
rect 660 462 716 478
rect 746 648 802 672
rect 746 614 757 648
rect 791 614 802 648
rect 746 580 802 614
rect 746 546 757 580
rect 791 546 802 580
rect 746 512 802 546
rect 746 478 757 512
rect 791 478 802 512
rect 746 462 802 478
rect 832 648 888 672
rect 832 614 843 648
rect 877 614 888 648
rect 832 580 888 614
rect 832 546 843 580
rect 877 546 888 580
rect 832 512 888 546
rect 832 478 843 512
rect 877 478 888 512
rect 832 462 888 478
rect 918 648 974 672
rect 918 614 929 648
rect 963 614 974 648
rect 918 580 974 614
rect 918 546 929 580
rect 963 546 974 580
rect 918 512 974 546
rect 918 478 929 512
rect 963 478 974 512
rect 918 462 974 478
rect 1004 648 1057 672
rect 1004 614 1015 648
rect 1049 614 1057 648
rect 1004 580 1057 614
rect 1004 546 1015 580
rect 1049 546 1057 580
rect 1004 512 1057 546
rect 1004 478 1015 512
rect 1049 478 1057 512
rect 1004 462 1057 478
<< ndiffc >>
rect 155 1790 189 1824
rect 155 1722 189 1756
rect 155 1654 189 1688
rect 241 1790 275 1824
rect 241 1722 275 1756
rect 241 1654 275 1688
rect 327 1790 361 1824
rect 327 1722 361 1756
rect 327 1654 361 1688
rect 413 1790 447 1824
rect 413 1722 447 1756
rect 413 1654 447 1688
rect 499 1790 533 1824
rect 499 1722 533 1756
rect 499 1654 533 1688
rect 585 1790 619 1824
rect 585 1722 619 1756
rect 585 1654 619 1688
rect 671 1790 705 1824
rect 671 1722 705 1756
rect 671 1654 705 1688
rect 757 1790 791 1824
rect 757 1722 791 1756
rect 757 1654 791 1688
rect 843 1790 877 1824
rect 843 1722 877 1756
rect 843 1654 877 1688
rect 929 1790 963 1824
rect 929 1722 963 1756
rect 929 1654 963 1688
rect 1015 1790 1049 1824
rect 1015 1722 1049 1756
rect 1015 1654 1049 1688
rect 155 614 189 648
rect 155 546 189 580
rect 155 478 189 512
rect 241 614 275 648
rect 241 546 275 580
rect 241 478 275 512
rect 327 614 361 648
rect 327 546 361 580
rect 327 478 361 512
rect 413 614 447 648
rect 413 546 447 580
rect 413 478 447 512
rect 499 614 533 648
rect 499 546 533 580
rect 499 478 533 512
rect 585 614 619 648
rect 585 546 619 580
rect 585 478 619 512
rect 671 614 705 648
rect 671 546 705 580
rect 671 478 705 512
rect 757 614 791 648
rect 757 546 791 580
rect 757 478 791 512
rect 843 614 877 648
rect 843 546 877 580
rect 843 478 877 512
rect 929 614 963 648
rect 929 546 963 580
rect 929 478 963 512
rect 1015 614 1049 648
rect 1015 546 1049 580
rect 1015 478 1049 512
<< psubdiff >>
rect 241 2537 275 2632
rect 241 2408 275 2503
rect 413 2537 447 2632
rect 413 2408 447 2503
rect 585 2537 619 2632
rect 585 2408 619 2503
rect 757 2537 791 2632
rect 757 2408 791 2503
rect 929 2537 963 2632
rect 929 2408 963 2503
<< psubdiffcont >>
rect 241 2503 275 2537
rect 413 2503 447 2537
rect 585 2503 619 2537
rect 757 2503 791 2537
rect 929 2503 963 2537
<< poly >>
rect 200 2117 316 2127
rect 200 2083 241 2117
rect 275 2083 316 2117
rect 200 2073 316 2083
rect 200 1848 230 2073
rect 286 1848 316 2073
rect 372 2117 488 2127
rect 372 2083 413 2117
rect 447 2083 488 2117
rect 372 2073 488 2083
rect 372 1848 402 2073
rect 458 1848 488 2073
rect 544 2117 660 2127
rect 544 2083 585 2117
rect 619 2083 660 2117
rect 544 2073 660 2083
rect 544 1848 574 2073
rect 630 1848 660 2073
rect 716 2117 832 2127
rect 716 2083 757 2117
rect 791 2083 832 2117
rect 716 2073 832 2083
rect 716 1848 746 2073
rect 802 1848 832 2073
rect 888 2117 1004 2127
rect 888 2083 929 2117
rect 963 2083 1004 2117
rect 888 2073 1004 2083
rect 888 1848 918 2073
rect 974 1848 1004 2073
rect 200 1428 230 1638
rect 286 1428 316 1638
rect 372 1428 402 1638
rect 458 1428 488 1638
rect 544 1428 574 1638
rect 630 1428 660 1638
rect 716 1428 746 1638
rect 802 1428 832 1638
rect 888 1428 918 1638
rect 974 1428 1004 1638
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 672 230 897
rect 286 672 316 897
rect 372 941 488 951
rect 372 907 413 941
rect 447 907 488 941
rect 372 897 488 907
rect 372 672 402 897
rect 458 672 488 897
rect 544 941 660 951
rect 544 907 585 941
rect 619 907 660 941
rect 544 897 660 907
rect 544 672 574 897
rect 630 672 660 897
rect 716 941 832 951
rect 716 907 757 941
rect 791 907 832 941
rect 716 897 832 907
rect 716 672 746 897
rect 802 672 832 897
rect 888 941 1004 951
rect 888 907 929 941
rect 963 907 1004 941
rect 888 897 1004 907
rect 888 672 918 897
rect 974 672 1004 897
rect 200 252 230 462
rect 286 252 316 462
rect 372 252 402 462
rect 458 252 488 462
rect 544 252 574 462
rect 630 252 660 462
rect 716 252 746 462
rect 802 252 832 462
rect 888 252 918 462
rect 974 252 1004 462
<< polycont >>
rect 241 2083 275 2117
rect 413 2083 447 2117
rect 585 2083 619 2117
rect 757 2083 791 2117
rect 929 2083 963 2117
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
<< locali >>
rect 233 2537 283 2621
rect 233 2503 241 2537
rect 275 2503 283 2537
rect 233 2419 283 2503
rect 405 2537 455 2621
rect 405 2503 413 2537
rect 447 2503 455 2537
rect 405 2419 455 2503
rect 577 2537 627 2621
rect 577 2503 585 2537
rect 619 2503 627 2537
rect 577 2419 627 2503
rect 749 2537 799 2621
rect 749 2503 757 2537
rect 791 2503 799 2537
rect 749 2419 799 2503
rect 921 2537 971 2621
rect 921 2503 929 2537
rect 963 2503 971 2537
rect 921 2419 971 2503
rect 233 2117 283 2201
rect 233 2083 241 2117
rect 275 2083 283 2117
rect 233 1999 283 2083
rect 405 2117 455 2201
rect 405 2083 413 2117
rect 447 2083 455 2117
rect 405 1999 455 2083
rect 577 2117 627 2201
rect 577 2083 585 2117
rect 619 2083 627 2117
rect 577 1999 627 2083
rect 749 2117 799 2201
rect 749 2083 757 2117
rect 791 2083 799 2117
rect 749 1999 799 2083
rect 921 2117 971 2201
rect 921 2083 929 2117
rect 963 2083 971 2117
rect 921 1999 971 2083
rect 147 1824 197 1949
rect 147 1790 155 1824
rect 189 1790 197 1824
rect 147 1756 197 1790
rect 147 1722 155 1756
rect 189 1722 197 1756
rect 147 1688 197 1722
rect 147 1654 155 1688
rect 189 1654 197 1688
rect 147 1361 197 1654
rect 147 1327 155 1361
rect 189 1327 197 1361
rect 147 1243 197 1327
rect 233 1824 283 1949
rect 233 1790 241 1824
rect 275 1790 283 1824
rect 233 1756 283 1790
rect 233 1722 241 1756
rect 275 1722 283 1756
rect 233 1688 283 1722
rect 233 1654 241 1688
rect 275 1654 283 1688
rect 233 1277 283 1654
rect 233 1243 241 1277
rect 275 1243 283 1277
rect 319 1824 369 1949
rect 319 1790 327 1824
rect 361 1790 369 1824
rect 319 1756 369 1790
rect 319 1722 327 1756
rect 361 1722 369 1756
rect 319 1688 369 1722
rect 319 1654 327 1688
rect 361 1654 369 1688
rect 319 1361 369 1654
rect 319 1327 327 1361
rect 361 1327 369 1361
rect 319 1243 369 1327
rect 405 1824 455 1949
rect 405 1790 413 1824
rect 447 1790 455 1824
rect 405 1756 455 1790
rect 405 1722 413 1756
rect 447 1722 455 1756
rect 405 1688 455 1722
rect 405 1654 413 1688
rect 447 1654 455 1688
rect 405 1277 455 1654
rect 405 1243 413 1277
rect 447 1243 455 1277
rect 491 1824 541 1949
rect 491 1790 499 1824
rect 533 1790 541 1824
rect 491 1756 541 1790
rect 491 1722 499 1756
rect 533 1722 541 1756
rect 491 1688 541 1722
rect 491 1654 499 1688
rect 533 1654 541 1688
rect 491 1361 541 1654
rect 491 1327 499 1361
rect 533 1327 541 1361
rect 491 1243 541 1327
rect 577 1824 627 1949
rect 577 1790 585 1824
rect 619 1790 627 1824
rect 577 1756 627 1790
rect 577 1722 585 1756
rect 619 1722 627 1756
rect 577 1688 627 1722
rect 577 1654 585 1688
rect 619 1654 627 1688
rect 577 1277 627 1654
rect 577 1243 585 1277
rect 619 1243 627 1277
rect 663 1824 713 1949
rect 663 1790 671 1824
rect 705 1790 713 1824
rect 663 1756 713 1790
rect 663 1722 671 1756
rect 705 1722 713 1756
rect 663 1688 713 1722
rect 663 1654 671 1688
rect 705 1654 713 1688
rect 663 1361 713 1654
rect 663 1327 671 1361
rect 705 1327 713 1361
rect 663 1243 713 1327
rect 749 1824 799 1949
rect 749 1790 757 1824
rect 791 1790 799 1824
rect 749 1756 799 1790
rect 749 1722 757 1756
rect 791 1722 799 1756
rect 749 1688 799 1722
rect 749 1654 757 1688
rect 791 1654 799 1688
rect 749 1277 799 1654
rect 749 1243 757 1277
rect 791 1243 799 1277
rect 835 1824 885 1949
rect 835 1790 843 1824
rect 877 1790 885 1824
rect 835 1756 885 1790
rect 835 1722 843 1756
rect 877 1722 885 1756
rect 835 1688 885 1722
rect 835 1654 843 1688
rect 877 1654 885 1688
rect 835 1361 885 1654
rect 835 1327 843 1361
rect 877 1327 885 1361
rect 835 1243 885 1327
rect 921 1824 971 1949
rect 921 1790 929 1824
rect 963 1790 971 1824
rect 921 1756 971 1790
rect 921 1722 929 1756
rect 963 1722 971 1756
rect 921 1688 971 1722
rect 921 1654 929 1688
rect 963 1654 971 1688
rect 921 1277 971 1654
rect 921 1243 929 1277
rect 963 1243 971 1277
rect 1007 1824 1057 1949
rect 1007 1790 1015 1824
rect 1049 1790 1057 1824
rect 1007 1756 1057 1790
rect 1007 1722 1015 1756
rect 1049 1722 1057 1756
rect 1007 1688 1057 1722
rect 1007 1654 1015 1688
rect 1049 1654 1057 1688
rect 1007 1361 1057 1654
rect 1007 1327 1015 1361
rect 1049 1327 1057 1361
rect 1007 1243 1057 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 405 941 455 1025
rect 405 907 413 941
rect 447 907 455 941
rect 405 823 455 907
rect 577 941 627 1025
rect 577 907 585 941
rect 619 907 627 941
rect 577 823 627 907
rect 749 941 799 1025
rect 749 907 757 941
rect 791 907 799 941
rect 749 823 799 907
rect 921 941 971 1025
rect 921 907 929 941
rect 963 907 971 941
rect 921 823 971 907
rect 147 648 197 773
rect 147 614 155 648
rect 189 614 197 648
rect 147 580 197 614
rect 147 546 155 580
rect 189 546 197 580
rect 147 512 197 546
rect 147 478 155 512
rect 189 478 197 512
rect 147 185 197 478
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 648 283 773
rect 233 614 241 648
rect 275 614 283 648
rect 233 580 283 614
rect 233 546 241 580
rect 275 546 283 580
rect 233 512 283 546
rect 233 478 241 512
rect 275 478 283 512
rect 233 101 283 478
rect 233 67 241 101
rect 275 67 283 101
rect 319 648 369 773
rect 319 614 327 648
rect 361 614 369 648
rect 319 580 369 614
rect 319 546 327 580
rect 361 546 369 580
rect 319 512 369 546
rect 319 478 327 512
rect 361 478 369 512
rect 319 185 369 478
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
rect 405 648 455 773
rect 405 614 413 648
rect 447 614 455 648
rect 405 580 455 614
rect 405 546 413 580
rect 447 546 455 580
rect 405 512 455 546
rect 405 478 413 512
rect 447 478 455 512
rect 405 101 455 478
rect 405 67 413 101
rect 447 67 455 101
rect 491 648 541 773
rect 491 614 499 648
rect 533 614 541 648
rect 491 580 541 614
rect 491 546 499 580
rect 533 546 541 580
rect 491 512 541 546
rect 491 478 499 512
rect 533 478 541 512
rect 491 185 541 478
rect 491 151 499 185
rect 533 151 541 185
rect 491 67 541 151
rect 577 648 627 773
rect 577 614 585 648
rect 619 614 627 648
rect 577 580 627 614
rect 577 546 585 580
rect 619 546 627 580
rect 577 512 627 546
rect 577 478 585 512
rect 619 478 627 512
rect 577 101 627 478
rect 577 67 585 101
rect 619 67 627 101
rect 663 648 713 773
rect 663 614 671 648
rect 705 614 713 648
rect 663 580 713 614
rect 663 546 671 580
rect 705 546 713 580
rect 663 512 713 546
rect 663 478 671 512
rect 705 478 713 512
rect 663 185 713 478
rect 663 151 671 185
rect 705 151 713 185
rect 663 67 713 151
rect 749 648 799 773
rect 749 614 757 648
rect 791 614 799 648
rect 749 580 799 614
rect 749 546 757 580
rect 791 546 799 580
rect 749 512 799 546
rect 749 478 757 512
rect 791 478 799 512
rect 749 101 799 478
rect 749 67 757 101
rect 791 67 799 101
rect 835 648 885 773
rect 835 614 843 648
rect 877 614 885 648
rect 835 580 885 614
rect 835 546 843 580
rect 877 546 885 580
rect 835 512 885 546
rect 835 478 843 512
rect 877 478 885 512
rect 835 185 885 478
rect 835 151 843 185
rect 877 151 885 185
rect 835 67 885 151
rect 921 648 971 773
rect 921 614 929 648
rect 963 614 971 648
rect 921 580 971 614
rect 921 546 929 580
rect 963 546 971 580
rect 921 512 971 546
rect 921 478 929 512
rect 963 478 971 512
rect 921 101 971 478
rect 921 67 929 101
rect 963 67 971 101
rect 1007 648 1057 773
rect 1007 614 1015 648
rect 1049 614 1057 648
rect 1007 580 1057 614
rect 1007 546 1015 580
rect 1049 546 1057 580
rect 1007 512 1057 546
rect 1007 478 1015 512
rect 1049 478 1057 512
rect 1007 185 1057 478
rect 1007 151 1015 185
rect 1049 151 1057 185
rect 1007 67 1057 151
<< viali >>
rect 241 2503 275 2537
rect 413 2503 447 2537
rect 585 2503 619 2537
rect 757 2503 791 2537
rect 929 2503 963 2537
rect 241 2083 275 2117
rect 413 2083 447 2117
rect 585 2083 619 2117
rect 757 2083 791 2117
rect 929 2083 963 2117
rect 155 1327 189 1361
rect 241 1243 275 1277
rect 327 1327 361 1361
rect 413 1243 447 1277
rect 499 1327 533 1361
rect 585 1243 619 1277
rect 671 1327 705 1361
rect 757 1243 791 1277
rect 843 1327 877 1361
rect 929 1243 963 1277
rect 1015 1327 1049 1361
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
rect 413 67 447 101
rect 499 151 533 185
rect 585 67 619 101
rect 671 151 705 185
rect 757 67 791 101
rect 843 151 877 185
rect 929 67 963 101
rect 1015 151 1049 185
<< metal1 >>
rect 224 2546 980 2548
rect 224 2537 662 2546
rect 224 2503 241 2537
rect 275 2503 413 2537
rect 447 2503 585 2537
rect 619 2503 662 2537
rect 224 2494 662 2503
rect 714 2537 980 2546
rect 714 2503 757 2537
rect 791 2503 929 2537
rect 963 2503 980 2537
rect 714 2494 980 2503
rect 224 2492 980 2494
rect 224 2126 980 2128
rect 224 2117 576 2126
rect 628 2117 980 2126
rect 224 2083 241 2117
rect 275 2083 413 2117
rect 447 2083 576 2117
rect 628 2083 757 2117
rect 791 2083 929 2117
rect 963 2083 980 2117
rect 224 2074 576 2083
rect 628 2074 980 2083
rect 224 2072 980 2074
rect 138 1370 1066 1372
rect 138 1361 662 1370
rect 714 1361 1066 1370
rect 138 1327 155 1361
rect 189 1327 327 1361
rect 361 1327 499 1361
rect 533 1327 662 1361
rect 714 1327 843 1361
rect 877 1327 1015 1361
rect 1049 1327 1066 1361
rect 138 1318 662 1327
rect 714 1318 1066 1327
rect 138 1316 1066 1318
rect 224 1286 980 1288
rect 224 1277 490 1286
rect 224 1243 241 1277
rect 275 1243 413 1277
rect 447 1243 490 1277
rect 224 1234 490 1243
rect 542 1277 980 1286
rect 542 1243 585 1277
rect 619 1243 757 1277
rect 791 1243 929 1277
rect 963 1243 980 1277
rect 542 1234 980 1243
rect 224 1232 980 1234
rect 224 950 980 952
rect 224 941 576 950
rect 628 941 980 950
rect 224 907 241 941
rect 275 907 413 941
rect 447 907 576 941
rect 628 907 757 941
rect 791 907 929 941
rect 963 907 980 941
rect 224 898 576 907
rect 628 898 980 907
rect 224 896 980 898
rect 138 194 1066 196
rect 138 185 662 194
rect 714 185 1066 194
rect 138 151 155 185
rect 189 151 327 185
rect 361 151 499 185
rect 533 151 662 185
rect 714 151 843 185
rect 877 151 1015 185
rect 1049 151 1066 185
rect 138 142 662 151
rect 714 142 1066 151
rect 138 140 1066 142
rect 224 110 980 112
rect 224 101 490 110
rect 224 67 241 101
rect 275 67 413 101
rect 447 67 490 101
rect 224 58 490 67
rect 542 101 980 110
rect 542 67 585 101
rect 619 67 757 101
rect 791 67 929 101
rect 963 67 980 101
rect 542 58 980 67
rect 224 56 980 58
<< via1 >>
rect 662 2494 714 2546
rect 576 2117 628 2126
rect 576 2083 585 2117
rect 585 2083 619 2117
rect 619 2083 628 2117
rect 576 2074 628 2083
rect 662 1361 714 1370
rect 662 1327 671 1361
rect 671 1327 705 1361
rect 705 1327 714 1361
rect 662 1318 714 1327
rect 490 1234 542 1286
rect 576 941 628 950
rect 576 907 585 941
rect 585 907 619 941
rect 619 907 628 941
rect 576 898 628 907
rect 662 185 714 194
rect 662 151 671 185
rect 671 151 705 185
rect 705 151 714 185
rect 662 142 714 151
rect 490 58 542 110
<< metal2 >>
rect 660 2546 716 2552
rect 660 2494 662 2546
rect 714 2494 716 2546
rect 574 2126 630 2132
rect 574 2074 576 2126
rect 628 2074 630 2126
rect 488 1286 544 1292
rect 488 1234 490 1286
rect 542 1234 544 1286
rect 488 110 544 1234
rect 574 950 630 2074
rect 574 898 576 950
rect 628 898 630 950
rect 574 892 630 898
rect 660 1370 716 2494
rect 660 1318 662 1370
rect 714 1318 716 1370
rect 660 194 716 1318
rect 660 142 662 194
rect 714 142 716 194
rect 660 136 716 142
rect 488 58 490 110
rect 542 58 544 110
rect 488 52 544 58
<< end >>
