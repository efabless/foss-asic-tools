magic
tech sky130A
magscale 1 2
timestamp 1621838304
<< xpolycontact >>
rect -141 2000 141 2432
rect -141 -2432 141 -2000
<< ppolyres >>
rect -141 -2000 141 2000
<< viali >>
rect -125 2017 125 2414
rect -125 -2414 125 -2017
<< metal1 >>
rect -131 2414 131 2426
rect -131 2017 -125 2414
rect 125 2017 131 2414
rect -131 2005 131 2017
rect -131 -2017 131 -2005
rect -131 -2414 -125 -2017
rect 125 -2414 131 -2017
rect -131 -2426 131 -2414
<< res1p41 >>
rect -143 -2002 143 2002
<< properties >>
string gencell sky130_fd_pr__res_high_po_1p41
string parameters w 1.410 l 20 m 1 nx 1 wmin 1.410 lmin 0.50 rho 319.8 val 4.563k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
