magic
tech sky130A
magscale 1 2
timestamp 1621758535
<< xpolycontact >>
rect -141 3000 141 3432
rect -141 -3432 141 -3000
<< ppolyres >>
rect -141 -3000 141 3000
<< viali >>
rect -125 3017 125 3414
rect -125 -3414 125 -3017
<< metal1 >>
rect -131 3414 131 3426
rect -131 3017 -125 3414
rect 125 3017 131 3414
rect -131 3005 131 3017
rect -131 -3017 131 -3005
rect -131 -3414 -125 -3017
rect 125 -3414 131 -3017
rect -131 -3426 131 -3414
<< res1p41 >>
rect -143 -3002 143 3002
<< properties >>
string gencell sky130_fd_pr__res_high_po_1p41
string parameters w 1.410 l 30 m 1 nx 1 wmin 1.410 lmin 0.50 rho 319.8 val 6.831k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
