magic
tech sky130A
magscale 1 2
timestamp 1622253817
<< nwell >>
rect -9000 40 9000 4500
<< pwell >>
rect -9000 -4500 9000 -40
<< mvpsubdiff >>
rect -8934 -118 8934 -106
rect -8934 -278 -8700 -118
rect 8700 -278 8934 -118
rect -8934 -290 8934 -278
rect -8934 -340 -8750 -290
rect -8934 -4200 -8922 -340
rect -8762 -4200 -8750 -340
rect -8934 -4250 -8750 -4200
rect 8750 -340 8934 -290
rect 8750 -4200 8762 -340
rect 8922 -4200 8934 -340
rect 8750 -4250 8934 -4200
rect -8934 -4262 8934 -4250
rect -8934 -4422 -8700 -4262
rect 8700 -4422 8934 -4262
rect -8934 -4434 8934 -4422
<< mvnsubdiff >>
rect -8934 4422 8934 4434
rect -8934 4262 -8700 4422
rect 8700 4262 8934 4422
rect -8934 4250 8934 4262
rect -8934 4200 -8750 4250
rect -8934 340 -8922 4200
rect -8762 340 -8750 4200
rect -8934 290 -8750 340
rect 8750 4200 8934 4250
rect 8750 340 8762 4200
rect 8922 340 8934 4200
rect 8750 290 8934 340
rect -8934 278 8934 290
rect -8934 118 -8700 278
rect 8700 118 8934 278
rect -8934 106 8934 118
<< mvpsubdiffcont >>
rect -8700 -278 8700 -118
rect -8922 -4200 -8762 -340
rect 8762 -4200 8922 -340
rect -8700 -4422 8700 -4262
<< mvnsubdiffcont >>
rect -8700 4262 8700 4422
rect -8922 340 -8762 4200
rect 8762 340 8922 4200
rect -8700 118 8700 278
<< locali >>
rect -8922 4200 -8762 4422
rect 8762 4200 8922 4422
rect 236 2511 336 2512
rect -1743 2502 1743 2511
rect -1743 2444 255 2502
rect 313 2444 1743 2502
rect -1743 2232 1743 2444
rect -1743 2172 -1611 2232
rect -1485 2172 -1353 2232
rect -711 2172 -579 2232
rect -453 2172 -321 2232
rect 321 2172 453 2232
rect 579 2172 711 2232
rect 1353 2172 1485 2232
rect 1611 2172 1743 2232
rect -4323 979 -4191 1028
rect -3807 979 -3675 1028
rect -3291 992 -3159 1028
rect -3033 992 -2901 1028
rect -2775 992 -2643 1028
rect -2517 992 -2385 1028
rect -2259 992 -2127 1028
rect -2001 992 -1869 1028
rect -3291 979 -1869 992
rect -1227 992 -1095 1028
rect -969 992 -837 1028
rect -1227 979 -837 992
rect -195 992 -63 1028
rect 63 992 195 1028
rect -195 979 195 992
rect 837 992 969 1028
rect 1095 992 1227 1028
rect 837 979 1227 992
rect 1869 992 2001 1028
rect 2127 992 2259 1028
rect 2385 992 2517 1028
rect 2643 992 2775 1028
rect 2901 992 3033 1028
rect 3159 992 3291 1028
rect 1869 979 3291 992
rect 3675 979 3807 1028
rect 4191 979 4323 1028
rect -4323 958 4323 979
rect -4323 949 -27 958
rect 29 949 4323 958
rect -4323 891 -28 949
rect 32 891 4323 949
rect -4323 823 4323 891
rect -8922 118 -8762 340
rect 8762 118 8922 340
rect -8922 -340 -8762 -118
rect 8762 -340 8922 -118
rect -4839 -3784 -1353 -3547
rect -4839 -3842 -2349 -3784
rect -2291 -3842 -1353 -3784
rect -4839 -3868 -1353 -3842
rect -8922 -4422 -8762 -4200
rect 8762 -4422 8922 -4200
<< viali >>
rect -8762 4262 -8700 4422
rect -8700 4262 8700 4422
rect 8700 4262 8762 4422
rect -8922 477 -8762 4063
rect 255 2444 313 2502
rect -27 949 29 958
rect -28 891 32 949
rect 8762 477 8922 4063
rect -8762 118 -8700 278
rect -8700 118 8700 278
rect 8700 118 8762 278
rect -8762 -278 -8700 -118
rect -8700 -278 8700 -118
rect 8700 -278 8762 -118
rect -8922 -4063 -8762 -477
rect -2349 -3842 -2291 -3784
rect 8762 -4063 8922 -477
rect -8762 -4422 -8700 -4262
rect -8700 -4422 8700 -4262
rect 8700 -4422 8762 -4262
<< metal1 >>
rect -8928 4422 8928 4428
rect -8928 4262 -8762 4422
rect 8762 4262 8928 4422
rect -8928 4256 8928 4262
rect -8928 4063 -8756 4256
rect -8928 477 -8922 4063
rect -8762 477 -8756 4063
rect -8156 3956 -8146 4256
rect -4667 2328 -4567 4256
rect -2372 2328 -2272 4256
rect -50 2328 50 4256
rect 243 2502 325 2508
rect 243 2444 255 2502
rect 313 2444 325 2502
rect 243 2438 325 2444
rect 2272 2328 2372 4256
rect 4567 2328 4667 4256
rect 8146 3956 8156 4256
rect 8756 4063 8928 4256
rect -4667 2228 4667 2328
rect -4667 2100 -4621 2228
rect -4561 2178 -4469 2228
rect -4425 2130 -4415 2188
rect -4357 2130 -4211 2188
rect -4409 2100 -4363 2130
rect -4151 2100 -4105 2228
rect -4045 2178 -3953 2228
rect -3635 2100 -3589 2228
rect -3529 2178 -3437 2228
rect -3119 2100 -3073 2228
rect -2603 2100 -2557 2228
rect -2087 2100 -2041 2228
rect -1055 2100 -1009 2228
rect -23 2100 23 2228
rect 1009 2100 1055 2228
rect 2041 2100 2087 2228
rect 2557 2100 2603 2228
rect 3073 2100 3119 2228
rect 3437 2178 3529 2228
rect 3589 2100 3635 2228
rect 3953 2178 4045 2228
rect 4105 2100 4151 2228
rect 4211 2130 4357 2188
rect 4415 2130 4425 2188
rect 4469 2178 4561 2228
rect 4363 2100 4409 2130
rect 4621 2100 4667 2228
rect -3893 764 -3847 1100
rect -3377 1000 -3331 1100
rect -3393 942 -3383 1000
rect -3325 942 -3315 1000
rect -2861 764 -2815 1100
rect -2345 1000 -2299 1100
rect -2361 942 -2351 1000
rect -2293 942 -2283 1000
rect -1829 764 -1783 1100
rect -3909 706 -3899 764
rect -3841 706 -3831 764
rect -2877 706 -2867 764
rect -2809 706 -2799 764
rect -1845 706 -1835 764
rect -1777 706 -1767 764
rect -1571 646 -1525 1100
rect -1313 764 -1267 1100
rect -797 1000 -751 1100
rect -813 942 -803 1000
rect -745 942 -735 1000
rect -539 882 -493 1100
rect -281 1000 -235 1100
rect -298 942 -287 1000
rect -229 942 -218 1000
rect -33 967 35 970
rect -555 824 -545 882
rect -487 824 -477 882
rect -1329 706 -1319 764
rect -1261 706 -1251 764
rect -1587 588 -1577 646
rect -1519 588 -1509 646
rect -8928 284 -8756 477
rect -298 378 -218 942
rect -298 320 -287 378
rect -229 320 -218 378
rect -40 958 40 967
rect -40 949 -27 958
rect 29 949 40 958
rect -40 891 -28 949
rect 32 891 40 949
rect -40 378 40 891
rect 235 764 281 1100
rect -40 320 -29 378
rect 29 320 40 378
rect 218 706 229 764
rect 287 706 298 764
rect 218 460 298 706
rect 493 646 539 1100
rect 605 825 616 883
rect 674 825 685 883
rect 605 646 685 825
rect 751 764 797 1100
rect 1267 1000 1313 1100
rect 1251 942 1261 1000
rect 1319 942 1329 1000
rect 1525 882 1571 1100
rect 1783 1000 1829 1100
rect 1767 942 1777 1000
rect 1835 942 1845 1000
rect 1509 824 1519 882
rect 1577 824 1587 882
rect 2299 764 2345 1100
rect 2815 1000 2861 1100
rect 2799 942 2809 1000
rect 2867 942 2877 1000
rect 3331 764 3377 1100
rect 3847 1000 3893 1100
rect 3831 942 3841 1000
rect 3899 942 3909 1000
rect 735 706 745 764
rect 803 706 813 764
rect 2283 706 2293 764
rect 2351 706 2361 764
rect 3315 706 3325 764
rect 3383 706 3393 764
rect 477 588 487 646
rect 545 588 555 646
rect 605 588 616 646
rect 674 588 685 646
rect 605 578 685 588
rect 8756 477 8762 4063
rect 8922 477 8928 4063
rect 218 378 297 460
rect 218 320 229 378
rect 287 320 297 378
rect 8756 284 8928 477
rect -8928 278 8928 284
rect -8928 118 -8762 278
rect 8762 118 8928 278
rect -8928 112 8928 118
rect -8928 -118 8928 -112
rect -8928 -278 -8762 -118
rect 8762 -278 8928 -118
rect -8928 -284 8928 -278
rect -8928 -477 -8756 -284
rect -39 -401 -29 -343
rect 29 -401 39 -343
rect 219 -401 229 -343
rect 287 -401 297 -343
rect -8928 -4063 -8922 -477
rect -8762 -4063 -8756 -477
rect -6489 -560 -6479 -502
rect -6421 -560 -6411 -502
rect -5457 -560 -5447 -502
rect -5389 -560 -5379 -502
rect -4425 -560 -4415 -502
rect -4357 -560 -4347 -502
rect -6473 -800 -6427 -560
rect -5973 -700 -5963 -642
rect -5905 -700 -5895 -642
rect -5957 -800 -5911 -700
rect -5441 -800 -5395 -560
rect -4941 -700 -4931 -642
rect -4873 -700 -4863 -642
rect -4925 -800 -4879 -700
rect -4409 -800 -4363 -560
rect -3393 -561 -3383 -503
rect -3325 -561 -3315 -503
rect -2361 -560 -2351 -502
rect -2293 -560 -2283 -502
rect -1329 -560 -1319 -502
rect -1261 -560 -1251 -502
rect -297 -560 -287 -502
rect -229 -560 -219 -502
rect -3909 -700 -3899 -642
rect -3841 -700 -3831 -642
rect -3893 -800 -3847 -700
rect -3377 -801 -3331 -561
rect -2877 -700 -2867 -642
rect -2809 -700 -2799 -642
rect -2861 -800 -2815 -700
rect -2345 -800 -2299 -560
rect -1845 -700 -1835 -642
rect -1777 -700 -1767 -642
rect -1829 -800 -1783 -700
rect -1313 -800 -1267 -560
rect -813 -700 -803 -642
rect -745 -700 -735 -642
rect -797 -800 -751 -700
rect -281 -800 -235 -560
rect -23 -713 23 -401
rect 219 -642 297 -401
rect 8756 -477 8928 -284
rect 735 -561 745 -503
rect 803 -561 813 -503
rect 1767 -560 1777 -502
rect 1835 -560 1845 -502
rect 2799 -560 2809 -502
rect 2867 -560 2877 -502
rect 3831 -560 3841 -502
rect 3899 -560 3909 -502
rect 4863 -560 4873 -502
rect 4931 -560 4941 -502
rect 5895 -560 5905 -502
rect 5963 -560 5973 -502
rect 219 -700 229 -642
rect 287 -700 297 -642
rect -175 -759 175 -713
rect -23 -800 23 -759
rect 235 -800 281 -700
rect 751 -801 797 -561
rect 1251 -700 1261 -642
rect 1319 -700 1329 -642
rect 1267 -800 1313 -700
rect 1783 -800 1829 -560
rect 2283 -700 2293 -642
rect 2351 -700 2361 -642
rect 2299 -800 2345 -700
rect 2815 -800 2861 -560
rect 3315 -700 3325 -642
rect 3383 -700 3393 -642
rect 3331 -800 3377 -700
rect 3847 -800 3893 -560
rect 4347 -700 4357 -642
rect 4415 -700 4425 -642
rect 4363 -800 4409 -700
rect 4879 -800 4925 -560
rect 5379 -700 5389 -642
rect 5447 -700 5457 -642
rect 5395 -800 5441 -700
rect 5911 -800 5957 -560
rect 6411 -700 6421 -642
rect 6479 -700 6489 -642
rect 6427 -800 6473 -700
rect -6989 -1842 -6943 -1800
rect -6731 -1842 -6685 -1800
rect -6989 -1887 -6685 -1842
rect -6989 -2137 -6943 -1887
rect -6731 -2137 -6685 -1887
rect -6625 -1917 -6533 -1832
rect -6367 -1917 -6275 -1832
rect -6635 -1977 -6625 -1917
rect -6533 -1977 -6523 -1917
rect -6377 -1977 -6367 -1917
rect -6275 -1977 -6265 -1917
rect -6215 -2137 -6169 -1800
rect -6109 -2037 -6017 -1847
rect -5851 -2037 -5759 -1854
rect -6119 -2097 -6109 -2037
rect -6017 -2097 -6007 -2037
rect -5861 -2097 -5851 -2037
rect -5759 -2097 -5749 -2037
rect -5699 -2137 -5653 -1800
rect -5593 -1917 -5501 -1832
rect -5335 -1917 -5243 -1832
rect -5603 -1977 -5593 -1917
rect -5501 -1977 -5491 -1917
rect -5345 -1977 -5335 -1917
rect -5243 -1977 -5233 -1917
rect -5183 -2137 -5137 -1800
rect -5077 -2037 -4985 -1838
rect -4819 -2037 -4727 -1846
rect -5087 -2097 -5077 -2037
rect -4985 -2097 -4975 -2037
rect -4829 -2097 -4819 -2037
rect -4727 -2097 -4717 -2037
rect -4667 -2137 -4621 -1800
rect -4561 -1917 -4469 -1831
rect -4303 -1917 -4211 -1830
rect -4571 -1977 -4561 -1917
rect -4469 -1977 -4459 -1917
rect -4313 -1977 -4303 -1917
rect -4211 -1977 -4201 -1917
rect -4151 -2137 -4105 -1800
rect -4045 -2037 -3953 -1851
rect -3787 -2037 -3695 -1846
rect -4055 -2097 -4045 -2037
rect -3953 -2097 -3943 -2037
rect -3797 -2097 -3787 -2037
rect -3695 -2097 -3685 -2037
rect -3635 -2137 -3589 -1800
rect -3529 -1917 -3437 -1832
rect -3271 -1917 -3179 -1832
rect -3539 -1977 -3529 -1917
rect -3437 -1977 -3427 -1917
rect -3281 -1977 -3271 -1917
rect -3179 -1977 -3169 -1917
rect -3119 -2137 -3073 -1800
rect -3013 -2037 -2921 -1836
rect -2755 -2037 -2663 -1839
rect -3023 -2097 -3013 -2037
rect -2921 -2097 -2911 -2037
rect -2765 -2097 -2755 -2037
rect -2663 -2097 -2653 -2037
rect -2603 -2137 -2557 -1800
rect -2497 -1917 -2405 -1832
rect -2239 -1917 -2147 -1832
rect -2507 -1977 -2497 -1917
rect -2405 -1977 -2395 -1917
rect -2249 -1977 -2239 -1917
rect -2147 -1977 -2137 -1917
rect -2087 -2137 -2041 -1800
rect -1981 -2037 -1889 -1841
rect -1723 -2037 -1631 -1844
rect -1991 -2097 -1981 -2037
rect -1889 -2097 -1879 -2037
rect -1733 -2097 -1723 -2037
rect -1631 -2097 -1621 -2037
rect -1571 -2137 -1525 -1800
rect -1465 -1917 -1373 -1832
rect -1207 -1917 -1115 -1832
rect -1475 -1977 -1465 -1917
rect -1373 -1977 -1363 -1917
rect -1217 -1977 -1207 -1917
rect -1115 -1977 -1105 -1917
rect -1055 -2137 -1009 -1800
rect -949 -2037 -857 -1840
rect -691 -2037 -599 -1845
rect -959 -2097 -949 -2037
rect -857 -2097 -847 -2037
rect -701 -2097 -691 -2037
rect -599 -2097 -589 -2037
rect -539 -2137 -493 -1800
rect -433 -1917 -341 -1832
rect -443 -1977 -433 -1917
rect -341 -1977 -331 -1917
rect 341 -2037 433 -1860
rect 331 -2097 341 -2037
rect 433 -2097 443 -2037
rect 493 -2137 539 -1800
rect 599 -1917 691 -1832
rect 857 -1917 949 -1832
rect 589 -1977 599 -1917
rect 691 -1977 701 -1917
rect 847 -1977 857 -1917
rect 949 -1977 959 -1917
rect 1009 -2137 1055 -1800
rect 1115 -2037 1207 -1841
rect 1373 -2037 1465 -1843
rect 1105 -2097 1115 -2037
rect 1207 -2097 1217 -2037
rect 1363 -2097 1373 -2037
rect 1465 -2097 1475 -2037
rect 1525 -2137 1571 -1800
rect 1631 -1917 1723 -1832
rect 1889 -1917 1981 -1832
rect 1621 -1977 1631 -1917
rect 1723 -1977 1733 -1917
rect 1879 -1977 1889 -1917
rect 1981 -1977 1991 -1917
rect 2041 -2137 2087 -1800
rect 2147 -2037 2239 -1836
rect 2405 -2037 2497 -1838
rect 2137 -2097 2147 -2037
rect 2239 -2097 2249 -2037
rect 2395 -2097 2405 -2037
rect 2497 -2097 2507 -2037
rect 2557 -2137 2603 -1800
rect 2663 -1917 2755 -1831
rect 2921 -1917 3013 -1832
rect 2653 -1977 2663 -1917
rect 2755 -1977 2765 -1917
rect 2911 -1977 2921 -1917
rect 3013 -1977 3023 -1917
rect 3073 -2137 3119 -1800
rect 3179 -2037 3271 -1841
rect 3437 -2037 3529 -1844
rect 3169 -2097 3179 -2037
rect 3271 -2097 3281 -2037
rect 3427 -2097 3437 -2037
rect 3529 -2097 3539 -2037
rect 3589 -2137 3635 -1800
rect 3695 -1917 3787 -1832
rect 3953 -1917 4045 -1832
rect 3685 -1977 3695 -1917
rect 3787 -1977 3797 -1917
rect 3943 -1977 3953 -1917
rect 4045 -1977 4055 -1917
rect 4105 -2137 4151 -1800
rect 4211 -2037 4303 -1836
rect 4469 -2037 4561 -1839
rect 4201 -2097 4211 -2037
rect 4303 -2097 4313 -2037
rect 4459 -2097 4469 -2037
rect 4561 -2097 4571 -2037
rect 4621 -2137 4667 -1800
rect 4727 -1917 4819 -1832
rect 4985 -1917 5077 -1832
rect 4717 -1977 4727 -1917
rect 4819 -1977 4829 -1917
rect 4975 -1977 4985 -1917
rect 5077 -1977 5087 -1917
rect 5137 -2137 5183 -1800
rect 5243 -2037 5335 -1842
rect 5501 -2037 5593 -1844
rect 5233 -2097 5243 -2037
rect 5335 -2097 5345 -2037
rect 5491 -2097 5501 -2037
rect 5593 -2097 5603 -2037
rect 5653 -2137 5699 -1800
rect 5759 -1917 5851 -1832
rect 6017 -1917 6109 -1831
rect 5749 -1977 5759 -1917
rect 5851 -1977 5861 -1917
rect 6007 -1977 6017 -1917
rect 6109 -1977 6119 -1917
rect 6169 -2137 6215 -1800
rect 6685 -1841 6731 -1800
rect 6943 -1841 6989 -1800
rect 6275 -2037 6367 -1842
rect 6533 -2037 6625 -1850
rect 6685 -1886 6989 -1841
rect 6265 -2097 6275 -2037
rect 6367 -2097 6377 -2037
rect 6523 -2097 6533 -2037
rect 6625 -2097 6635 -2037
rect 6685 -2137 6731 -1886
rect 6943 -2137 6989 -1886
rect -6989 -2217 6989 -2137
rect -63 -2257 63 -2217
rect 7114 -2239 7125 -2181
rect 7183 -2239 7194 -2181
rect 7114 -2257 7194 -2239
rect -4409 -2373 63 -2257
rect 2405 -2317 7194 -2257
rect -4409 -2500 -4363 -2373
rect -3893 -2500 -3847 -2373
rect -3377 -2500 -3331 -2373
rect -2861 -2500 -2815 -2373
rect -2345 -2500 -2299 -2373
rect -1829 -2500 -1783 -2373
rect 2405 -2468 2497 -2317
rect 2799 -2435 2809 -2377
rect 2867 -2435 2877 -2377
rect 2815 -2500 2861 -2435
rect 3179 -2468 3271 -2317
rect 3437 -2468 3529 -2317
rect 3847 -2500 3893 -2317
rect 4211 -2468 4303 -2317
rect 4469 -2468 4561 -2317
rect 4863 -2435 4873 -2377
rect 4931 -2435 4941 -2377
rect 4879 -2500 4925 -2435
rect 5243 -2468 5335 -2317
rect 5501 -2468 5593 -2317
rect 5911 -2500 5957 -2317
rect 6275 -2468 6367 -2317
rect -5189 -3541 -5131 -3500
rect -5189 -3587 -4985 -3541
rect -8928 -4256 -8756 -4063
rect -8156 -4256 -8146 -3956
rect -5189 -4256 -5131 -3587
rect -4925 -3600 -4879 -3500
rect -4941 -3658 -4931 -3600
rect -4873 -3658 -4863 -3600
rect -4673 -4256 -4615 -3500
rect -4157 -4256 -4099 -3500
rect -3641 -4256 -3583 -3500
rect -3125 -4256 -3067 -3500
rect -2609 -4256 -2551 -3500
rect -2361 -3784 -2279 -3778
rect -2361 -3842 -2349 -3784
rect -2291 -3842 -2279 -3784
rect -2361 -3848 -2279 -3842
rect -2093 -4256 -2035 -3500
rect -1577 -4256 -1519 -3500
rect -1313 -3600 -1267 -3500
rect -1061 -3541 -1003 -3500
rect -1207 -3587 -1003 -3541
rect -1329 -3658 -1319 -3600
rect -1261 -3658 -1251 -3600
rect -1061 -4256 -1003 -3587
rect 2041 -3541 2087 -3500
rect 2299 -3541 2345 -3500
rect 2041 -3587 2345 -3541
rect 2041 -4256 2087 -3587
rect 2299 -4256 2345 -3587
rect 2557 -3620 2603 -3500
rect 2541 -3678 2551 -3620
rect 2609 -3678 2619 -3620
rect 2663 -3947 2755 -3561
rect 2921 -3947 3013 -3562
rect 3073 -3620 3119 -3500
rect 3057 -3678 3067 -3620
rect 3125 -3678 3135 -3620
rect 2653 -4007 2663 -3947
rect 2755 -4007 2765 -3947
rect 2911 -4007 2921 -3947
rect 3013 -4007 3023 -3947
rect 3331 -4256 3377 -3500
rect 3589 -3788 3635 -3500
rect 3573 -3846 3583 -3788
rect 3641 -3846 3651 -3788
rect 3695 -3947 3787 -3556
rect 3953 -3947 4045 -3554
rect 4105 -3788 4151 -3500
rect 4089 -3846 4099 -3788
rect 4157 -3846 4167 -3788
rect 3685 -4007 3695 -3947
rect 3787 -4007 3797 -3947
rect 3943 -4007 3953 -3947
rect 4045 -4007 4055 -3947
rect 4363 -4256 4409 -3500
rect 4621 -3620 4667 -3500
rect 4605 -3678 4615 -3620
rect 4673 -3678 4683 -3620
rect 4727 -3947 4819 -3554
rect 4985 -3947 5077 -3553
rect 5137 -3620 5183 -3500
rect 5121 -3678 5131 -3620
rect 5189 -3678 5199 -3620
rect 4717 -4007 4727 -3947
rect 4819 -4007 4829 -3947
rect 4975 -4007 4985 -3947
rect 5077 -4007 5087 -3947
rect 5395 -4256 5441 -3500
rect 5653 -3788 5699 -3500
rect 5638 -3846 5648 -3788
rect 5706 -3846 5716 -3788
rect 5759 -3947 5851 -3553
rect 6017 -3947 6109 -3554
rect 6169 -3788 6215 -3500
rect 6427 -3541 6473 -3500
rect 6685 -3541 6731 -3500
rect 6427 -3587 6731 -3541
rect 6153 -3846 6163 -3788
rect 6221 -3846 6231 -3788
rect 5749 -4007 5759 -3947
rect 5851 -4007 5861 -3947
rect 6007 -4007 6017 -3947
rect 6109 -4007 6119 -3947
rect 6427 -4256 6473 -3587
rect 6685 -4256 6731 -3587
rect 8146 -4256 8156 -3956
rect 8756 -4063 8762 -477
rect 8922 -4063 8928 -477
rect 8756 -4256 8928 -4063
rect -8928 -4262 8928 -4256
rect -8928 -4422 -8762 -4262
rect 8762 -4422 8928 -4262
rect -8928 -4428 8928 -4422
<< via1 >>
rect -8756 3956 -8156 4256
rect 255 2444 313 2502
rect 8156 3956 8756 4256
rect -4415 2130 -4357 2188
rect 4357 2130 4415 2188
rect -3383 942 -3325 1000
rect -2351 942 -2293 1000
rect -3899 706 -3841 764
rect -2867 706 -2809 764
rect -1835 706 -1777 764
rect -803 942 -745 1000
rect -287 942 -229 1000
rect -545 824 -487 882
rect -1319 706 -1261 764
rect -1577 588 -1519 646
rect -287 320 -229 378
rect -29 320 29 378
rect 229 706 287 764
rect 616 825 674 883
rect 1261 942 1319 1000
rect 1777 942 1835 1000
rect 1519 824 1577 882
rect 2809 942 2867 1000
rect 3841 942 3899 1000
rect 745 706 803 764
rect 2293 706 2351 764
rect 3325 706 3383 764
rect 487 588 545 646
rect 616 588 674 646
rect 229 320 287 378
rect -29 -401 29 -343
rect 229 -401 287 -343
rect -6479 -560 -6421 -502
rect -5447 -560 -5389 -502
rect -4415 -560 -4357 -502
rect -5963 -700 -5905 -642
rect -4931 -700 -4873 -642
rect -3383 -561 -3325 -503
rect -2351 -560 -2293 -502
rect -1319 -560 -1261 -502
rect -287 -560 -229 -502
rect -3899 -700 -3841 -642
rect -2867 -700 -2809 -642
rect -1835 -700 -1777 -642
rect -803 -700 -745 -642
rect 745 -561 803 -503
rect 1777 -560 1835 -502
rect 2809 -560 2867 -502
rect 3841 -560 3899 -502
rect 4873 -560 4931 -502
rect 5905 -560 5963 -502
rect 229 -700 287 -642
rect 1261 -700 1319 -642
rect 2293 -700 2351 -642
rect 3325 -700 3383 -642
rect 4357 -700 4415 -642
rect 5389 -700 5447 -642
rect 6421 -700 6479 -642
rect -6625 -1977 -6533 -1917
rect -6367 -1977 -6275 -1917
rect -6109 -2097 -6017 -2037
rect -5851 -2097 -5759 -2037
rect -5593 -1977 -5501 -1917
rect -5335 -1977 -5243 -1917
rect -5077 -2097 -4985 -2037
rect -4819 -2097 -4727 -2037
rect -4561 -1977 -4469 -1917
rect -4303 -1977 -4211 -1917
rect -4045 -2097 -3953 -2037
rect -3787 -2097 -3695 -2037
rect -3529 -1977 -3437 -1917
rect -3271 -1977 -3179 -1917
rect -3013 -2097 -2921 -2037
rect -2755 -2097 -2663 -2037
rect -2497 -1977 -2405 -1917
rect -2239 -1977 -2147 -1917
rect -1981 -2097 -1889 -2037
rect -1723 -2097 -1631 -2037
rect -1465 -1977 -1373 -1917
rect -1207 -1977 -1115 -1917
rect -949 -2097 -857 -2037
rect -691 -2097 -599 -2037
rect -433 -1977 -341 -1917
rect 341 -2097 433 -2037
rect 599 -1977 691 -1917
rect 857 -1977 949 -1917
rect 1115 -2097 1207 -2037
rect 1373 -2097 1465 -2037
rect 1631 -1977 1723 -1917
rect 1889 -1977 1981 -1917
rect 2147 -2097 2239 -2037
rect 2405 -2097 2497 -2037
rect 2663 -1977 2755 -1917
rect 2921 -1977 3013 -1917
rect 3179 -2097 3271 -2037
rect 3437 -2097 3529 -2037
rect 3695 -1977 3787 -1917
rect 3953 -1977 4045 -1917
rect 4211 -2097 4303 -2037
rect 4469 -2097 4561 -2037
rect 4727 -1977 4819 -1917
rect 4985 -1977 5077 -1917
rect 5243 -2097 5335 -2037
rect 5501 -2097 5593 -2037
rect 5759 -1977 5851 -1917
rect 6017 -1977 6109 -1917
rect 6275 -2097 6367 -2037
rect 6533 -2097 6625 -2037
rect 7125 -2239 7183 -2181
rect 2809 -2435 2867 -2377
rect 4873 -2435 4931 -2377
rect -8756 -4256 -8156 -3956
rect -4931 -3658 -4873 -3600
rect -2349 -3842 -2291 -3784
rect -1319 -3658 -1261 -3600
rect 2551 -3678 2609 -3620
rect 3067 -3678 3125 -3620
rect 2663 -4007 2755 -3947
rect 2921 -4007 3013 -3947
rect 3583 -3846 3641 -3788
rect 4099 -3846 4157 -3788
rect 3695 -4007 3787 -3947
rect 3953 -4007 4045 -3947
rect 4615 -3678 4673 -3620
rect 5131 -3678 5189 -3620
rect 4727 -4007 4819 -3947
rect 4985 -4007 5077 -3947
rect 5648 -3846 5706 -3788
rect 6163 -3846 6221 -3788
rect 5759 -4007 5851 -3947
rect 6017 -4007 6109 -3947
rect 8156 -4256 8756 -3956
<< metal2 >>
rect -8756 4256 -8156 4266
rect -8756 3946 -8156 3956
rect 8156 4256 8756 4266
rect 8156 3946 8756 3956
rect 255 2502 313 2512
rect -5828 2390 50 2490
rect 255 2434 313 2444
rect -5828 968 -5708 2390
rect -50 2328 50 2390
rect -4415 2228 4415 2328
rect -4415 2188 -4357 2228
rect -4415 2120 -4357 2130
rect 4357 2188 4415 2228
rect 4357 2120 4415 2130
rect -7751 848 -5708 968
rect -3383 1000 3899 1010
rect -3325 942 -2351 1000
rect -2293 942 -803 1000
rect -745 942 -287 1000
rect -229 942 1261 1000
rect 1319 942 1777 1000
rect 1835 942 2809 1000
rect 2867 942 3841 1000
rect -3383 932 3899 942
rect 616 892 674 893
rect -545 883 1577 892
rect -545 882 616 883
rect -7751 -3708 -7631 848
rect -487 825 616 882
rect 674 882 1577 883
rect 674 825 1519 882
rect -487 824 1519 825
rect -545 814 1577 824
rect -3899 764 3383 774
rect -3841 706 -2867 764
rect -2809 706 -1835 764
rect -1777 706 -1319 764
rect -1261 706 229 764
rect 287 706 745 764
rect 803 706 2293 764
rect 2351 706 3325 764
rect -3899 696 3383 706
rect -1577 646 545 656
rect -1519 588 487 646
rect -1577 578 545 588
rect 616 646 7475 656
rect 674 643 7475 646
rect 674 588 7377 643
rect 616 578 7377 588
rect -555 538 -477 578
rect -555 458 7194 538
rect -298 378 -218 388
rect -298 320 -287 378
rect -229 320 -218 378
rect -298 -492 -218 320
rect -29 378 29 392
rect -29 -343 29 320
rect -29 -411 29 -401
rect 218 378 298 389
rect 218 320 229 378
rect 287 320 298 378
rect 218 -343 298 320
rect 218 -401 229 -343
rect 287 -401 298 -343
rect 218 -411 298 -401
rect -6479 -502 5963 -492
rect -6421 -560 -5447 -502
rect -5389 -560 -4415 -502
rect -4357 -503 -2351 -502
rect -4357 -560 -3383 -503
rect -6479 -561 -3383 -560
rect -3325 -560 -2351 -503
rect -2293 -560 -1319 -502
rect -1261 -560 -287 -502
rect -229 -503 1777 -502
rect -229 -560 745 -503
rect -3325 -561 745 -560
rect 803 -560 1777 -503
rect 1835 -560 2809 -502
rect 2867 -560 3841 -502
rect 3899 -560 4873 -502
rect 4931 -560 5905 -502
rect 803 -561 5963 -560
rect -6479 -570 5963 -561
rect -3383 -571 -3325 -570
rect 745 -571 803 -570
rect -5963 -642 6479 -632
rect -5905 -700 -4931 -642
rect -4873 -700 -3899 -642
rect -3841 -700 -2867 -642
rect -2809 -700 -1835 -642
rect -1777 -700 -803 -642
rect -745 -700 229 -642
rect 287 -700 1261 -642
rect 1319 -700 2293 -642
rect 2351 -700 3325 -642
rect 3383 -700 4357 -642
rect 4415 -700 5389 -642
rect 5447 -700 6421 -642
rect -5963 -710 6479 -700
rect -6625 -1917 6109 -1907
rect -6533 -1977 -6367 -1917
rect -6275 -1977 -5593 -1917
rect -5501 -1977 -5335 -1917
rect -5243 -1977 -4561 -1917
rect -4469 -1977 -4303 -1917
rect -4211 -1977 -3529 -1917
rect -3437 -1977 -3271 -1917
rect -3179 -1977 -2497 -1917
rect -2405 -1977 -2239 -1917
rect -2147 -1977 -1465 -1917
rect -1373 -1977 -1207 -1917
rect -1115 -1977 -433 -1917
rect -341 -1977 599 -1917
rect 691 -1977 857 -1917
rect 949 -1977 1631 -1917
rect 1723 -1977 1889 -1917
rect 1981 -1977 2663 -1917
rect 2755 -1977 2921 -1917
rect 3013 -1977 3695 -1917
rect 3787 -1977 3953 -1917
rect 4045 -1977 4727 -1917
rect 4819 -1977 4985 -1917
rect 5077 -1977 5759 -1917
rect 5851 -1977 6017 -1917
rect -6625 -1987 6109 -1977
rect -6625 -1997 -6533 -1987
rect -6625 -2055 -6612 -1997
rect -6554 -2055 -6533 -1997
rect -6625 -2064 -6533 -2055
rect -6109 -2037 6625 -2027
rect -6612 -2065 -6554 -2064
rect -6017 -2097 -5851 -2037
rect -5759 -2097 -5077 -2037
rect -4985 -2097 -4819 -2037
rect -4727 -2097 -4045 -2037
rect -3953 -2097 -3787 -2037
rect -3695 -2097 -3013 -2037
rect -2921 -2097 -2755 -2037
rect -2663 -2097 -1981 -2037
rect -1889 -2097 -1723 -2037
rect -1631 -2097 -949 -2037
rect -857 -2097 -691 -2037
rect -599 -2097 341 -2037
rect 433 -2097 1115 -2037
rect 1207 -2097 1373 -2037
rect 1465 -2097 2147 -2037
rect 2239 -2097 2405 -2037
rect 2497 -2097 3179 -2037
rect 3271 -2097 3437 -2037
rect 3529 -2097 4211 -2037
rect 4303 -2097 4469 -2037
rect 4561 -2097 5243 -2037
rect 5335 -2097 5501 -2037
rect 5593 -2097 6275 -2037
rect 6367 -2097 6533 -2037
rect -6109 -2107 6625 -2097
rect -6109 -2165 -6094 -2107
rect -6036 -2165 -6017 -2107
rect -6109 -2184 -6017 -2165
rect 7114 -2181 7194 458
rect 7275 443 7377 578
rect 7275 433 7475 443
rect 7275 59 7354 433
rect 7114 -2239 7125 -2181
rect 7183 -2239 7194 -2181
rect 7114 -2257 7194 -2239
rect 7274 -2337 7354 59
rect 2809 -2377 7354 -2337
rect 2867 -2397 4873 -2377
rect 2809 -2445 2867 -2435
rect 4931 -2397 7354 -2377
rect 4873 -2445 4931 -2435
rect -4931 -3600 -1261 -3590
rect -4873 -3658 -1319 -3600
rect -4931 -3668 -1261 -3658
rect 2551 -3620 2609 -3610
rect -3159 -3708 -3033 -3668
rect 3067 -3620 3125 -3610
rect 2609 -3678 3067 -3628
rect 4615 -3620 4673 -3610
rect 3125 -3678 4615 -3628
rect 5131 -3620 5189 -3610
rect 4673 -3678 5131 -3628
rect 2551 -3688 5189 -3678
rect -7756 -3828 -3033 -3708
rect 6283 -3750 6292 -3665
rect 6377 -3750 6386 -3665
rect -2349 -3784 -2291 -3774
rect -2349 -3852 -2291 -3842
rect 3583 -3788 3641 -3778
rect 4099 -3788 4157 -3778
rect 3641 -3846 4099 -3796
rect 5648 -3788 5706 -3778
rect 4157 -3846 5648 -3796
rect 6163 -3788 6221 -3778
rect 5706 -3846 6163 -3796
rect 3583 -3856 6221 -3846
rect 6287 -3937 6384 -3750
rect -8756 -3956 -8156 -3946
rect 2663 -3947 6384 -3937
rect 2755 -4007 2921 -3947
rect 3013 -4007 3695 -3947
rect 3787 -4007 3953 -3947
rect 4045 -4007 4727 -3947
rect 4819 -4007 4985 -3947
rect 5077 -4007 5759 -3947
rect 5851 -4007 6017 -3947
rect 6109 -4007 6384 -3947
rect 2663 -4017 6384 -4007
rect 8156 -3956 8756 -3946
rect -8756 -4266 -8156 -4256
rect 8156 -4266 8756 -4256
<< via2 >>
rect -8756 3956 -8156 4256
rect 8156 3956 8756 4256
rect 255 2444 313 2502
rect -6612 -2055 -6554 -1997
rect -6094 -2165 -6036 -2107
rect 7377 443 7475 643
rect 6292 -3750 6377 -3665
rect -2349 -3842 -2291 -3784
rect -8756 -4256 -8156 -3956
rect 8156 -4256 8756 -3956
<< metal3 >>
rect -8766 4256 -8146 4261
rect -8766 3956 -8756 4256
rect -8156 3956 -8146 4256
rect -8766 3951 -8146 3956
rect 8146 4256 8766 4261
rect 8146 3956 8156 4256
rect 8756 3956 8766 4256
rect 8146 3951 8766 3956
rect 233 2502 8680 2526
rect 233 2444 255 2502
rect 313 2444 8680 2502
rect 233 2426 8680 2444
rect 8580 2187 8680 2426
rect 8580 2087 9459 2187
rect 7367 643 7485 648
rect 7367 443 7377 643
rect 7475 443 7945 643
rect 7367 438 7485 443
rect -8700 132 -7304 232
rect -8700 -241 -7867 -141
rect -7967 -2250 -7867 -241
rect -7404 -1992 -7304 132
rect 7745 111 7945 443
rect 7745 -89 14651 111
rect 7969 -580 9459 -480
rect -7404 -1997 -6544 -1992
rect -7404 -2055 -6612 -1997
rect -6554 -2055 -6544 -1997
rect -7404 -2092 -6544 -2055
rect -6359 -2107 -6026 -2102
rect -6359 -2165 -6094 -2107
rect -6036 -2165 -6026 -2107
rect -6359 -2202 -6026 -2165
rect -6359 -2250 -6259 -2202
rect -7967 -2350 -6259 -2250
rect 7969 -2467 8064 -580
rect 6807 -2562 8064 -2467
rect 8333 -824 9449 -734
rect -8683 -2849 -5706 -2649
rect -8766 -3956 -8146 -3951
rect -8766 -4256 -8756 -3956
rect -8156 -4256 -8146 -3956
rect -5906 -3982 -5706 -2849
rect 6807 -3605 6902 -2562
rect 8333 -2833 8433 -824
rect 6287 -3665 6902 -3605
rect 6287 -3750 6292 -3665
rect 6377 -3700 6902 -3665
rect 6985 -2933 8433 -2833
rect 8604 -2862 9365 -2742
rect 6377 -3750 6382 -3700
rect 6287 -3755 6382 -3750
rect -2362 -3784 3150 -3767
rect -2362 -3842 -2349 -3784
rect -2291 -3815 3150 -3784
rect 6985 -3815 7085 -2933
rect 8604 -3049 8724 -2862
rect 8094 -3169 8724 -3049
rect 8094 -3351 8294 -3169
rect -2291 -3842 7085 -3815
rect -2362 -3867 7085 -3842
rect 3052 -3915 7085 -3867
rect 7290 -3551 8294 -3351
rect 7290 -3982 7490 -3551
rect -5906 -4182 7490 -3982
rect 8146 -3956 8766 -3951
rect -8766 -4261 -8146 -4256
rect 8146 -4256 8156 -3956
rect 8756 -4256 8766 -3956
rect 8146 -4261 8766 -4256
<< via3 >>
rect -8756 3956 -8156 4256
rect 8156 3956 8756 4256
rect -8756 -4256 -8156 -3956
rect 8156 -4256 8756 -3956
<< metal4 >>
rect -9000 4256 9000 4500
rect -9000 3956 -8756 4256
rect -8156 3956 8156 4256
rect 8756 3956 9000 4256
rect -9000 3700 9000 3956
rect -9000 -3956 9000 -3700
rect -9000 -4256 -8756 -3956
rect -8156 -4256 8156 -3956
rect 8756 -4256 9000 -3956
rect -9000 -4500 9000 -4256
<< comment >>
rect -19 -122 18 187
rect -3111 -2248 -3087 -2071
rect 4375 -2140 4394 -1995
use cascode_bias  cascode_bias_0 folded_cascode_p_in/./../bias-circuit
timestamp 1622253817
transform 1 0 12000 0 1 0
box -3000 -4500 3000 4500
use sky130_fd_pr__nfet_g5v0d10v5_7QEKRB  xm4 ../bias-circuit
timestamp 1621758535
transform 1 0 4386 0 1 -3000
box -2351 -588 2351 588
use sky130_fd_pr__nfet_g5v0d10v5_CQE3UR  xm3 ./../folded_cascode_n_in
timestamp 1620706892
transform 1 0 -3096 0 1 -3000
box -2093 -588 2093 588
use sky130_fd_pr__nfet_g5v0d10v5_3REK67  xm2 ./../folded_cascode_n_in
timestamp 1620706892
transform 1 0 0 0 1 -1300
box -6995 -588 6995 588
use sky130_fd_pr__pfet_g5v0d10v5_QUEZLW  xm1 ./../folded_cascode_n_in
timestamp 1620706892
transform 1 0 0 0 1 1600
box -4739 -600 4739 600
<< labels >>
flabel metal4 -9000 3700 -9000 4500 3 FreeSans 480 0 0 0 vdd
port 5 e
flabel metal4 -9000 -4500 -9000 -3700 3 FreeSans 480 0 0 0 vss
port 6 e
flabel metal3 -8700 132 -8700 232 1 FreeSans 240 0 0 0 in_m
port 2 n
flabel metal3 -8700 -241 -8700 -141 1 FreeSans 240 0 0 0 in_p
port 3 n
flabel metal3 -8683 -2849 -8683 -2649 1 FreeSans 240 0 0 0 ibias
port 1 n
flabel metal3 14651 -89 14651 111 1 FreeSans 240 0 0 0 out
port 4 n
<< properties >>
string FIXED_BBOX -8842 -4342 8842 -198
<< end >>
