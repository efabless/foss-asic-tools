magic
tech sky130A
magscale 1 2
timestamp 1678192885
<< nwell >>
rect 0 1512 516 3024
<< pwell >>
rect 121 814 395 1076
rect 215 30 301 306
<< nmos >>
rect 200 840 230 1050
rect 286 840 316 1050
<< pmos >>
rect 200 1995 230 2163
rect 286 1995 316 2163
<< ndiff >>
rect 147 1034 200 1050
rect 147 1000 155 1034
rect 189 1000 200 1034
rect 147 966 200 1000
rect 147 932 155 966
rect 189 932 200 966
rect 147 898 200 932
rect 147 864 155 898
rect 189 864 200 898
rect 147 840 200 864
rect 230 1034 286 1050
rect 230 1000 241 1034
rect 275 1000 286 1034
rect 230 966 286 1000
rect 230 932 241 966
rect 275 932 286 966
rect 230 898 286 932
rect 230 864 241 898
rect 275 864 286 898
rect 230 840 286 864
rect 316 1034 369 1050
rect 316 1000 327 1034
rect 361 1000 369 1034
rect 316 966 369 1000
rect 316 932 327 966
rect 361 932 369 966
rect 316 898 369 932
rect 316 864 327 898
rect 361 864 369 898
rect 316 840 369 864
<< pdiff >>
rect 147 2113 200 2163
rect 147 2079 155 2113
rect 189 2079 200 2113
rect 147 2045 200 2079
rect 147 2011 155 2045
rect 189 2011 200 2045
rect 147 1995 200 2011
rect 230 2113 286 2163
rect 230 2079 241 2113
rect 275 2079 286 2113
rect 230 2045 286 2079
rect 230 2011 241 2045
rect 275 2011 286 2045
rect 230 1995 286 2011
rect 316 2113 369 2163
rect 316 2079 327 2113
rect 361 2079 369 2113
rect 316 2045 369 2079
rect 316 2011 327 2045
rect 361 2011 369 2045
rect 316 1995 369 2011
<< ndiffc >>
rect 155 1000 189 1034
rect 155 932 189 966
rect 155 864 189 898
rect 241 1000 275 1034
rect 241 932 275 966
rect 241 864 275 898
rect 327 1000 361 1034
rect 327 932 361 966
rect 327 864 361 898
<< pdiffc >>
rect 155 2079 189 2113
rect 155 2011 189 2045
rect 241 2079 275 2113
rect 241 2011 275 2045
rect 327 2079 361 2113
rect 327 2011 361 2045
<< psubdiff >>
rect 241 185 275 280
rect 241 56 275 151
<< nsubdiff >>
rect 241 2873 275 2968
rect 241 2744 275 2839
<< psubdiffcont >>
rect 241 151 275 185
<< nsubdiffcont >>
rect 241 2839 275 2873
<< poly >>
rect 200 2453 316 2463
rect 200 2419 241 2453
rect 275 2419 316 2453
rect 200 2409 316 2419
rect 200 2163 230 2409
rect 286 2163 316 2409
rect 200 1764 230 1995
rect 286 1764 316 1995
rect 200 1050 230 1260
rect 286 1050 316 1260
rect 200 615 230 840
rect 286 615 316 840
rect 200 605 316 615
rect 200 571 241 605
rect 275 571 316 605
rect 200 561 316 571
<< polycont >>
rect 241 2419 275 2453
rect 241 571 275 605
<< locali >>
rect 233 2873 283 2957
rect 233 2839 241 2873
rect 275 2839 283 2873
rect 233 2755 283 2839
rect 233 2453 283 2537
rect 233 2419 241 2453
rect 275 2419 283 2453
rect 233 2335 283 2419
rect 147 2113 197 2285
rect 147 2079 155 2113
rect 189 2079 197 2113
rect 147 2045 197 2079
rect 147 2011 155 2045
rect 189 2011 197 2045
rect 147 1697 197 2011
rect 147 1663 155 1697
rect 189 1663 197 1697
rect 147 1579 197 1663
rect 233 2113 283 2285
rect 233 2079 241 2113
rect 275 2079 283 2113
rect 233 2045 283 2079
rect 233 2011 241 2045
rect 275 2011 283 2045
rect 233 1613 283 2011
rect 233 1579 241 1613
rect 275 1579 283 1613
rect 319 2113 369 2285
rect 319 2079 327 2113
rect 361 2079 369 2113
rect 319 2045 369 2079
rect 319 2011 327 2045
rect 361 2011 369 2045
rect 319 1697 369 2011
rect 319 1663 327 1697
rect 361 1663 369 1697
rect 319 1579 369 1663
rect 405 1579 413 1613
rect 447 1579 455 1613
rect 405 1445 455 1579
rect 147 1361 197 1445
rect 147 1327 155 1361
rect 189 1327 197 1361
rect 147 1034 197 1327
rect 147 1000 155 1034
rect 189 1000 197 1034
rect 147 966 197 1000
rect 147 932 155 966
rect 189 932 197 966
rect 147 898 197 932
rect 147 864 155 898
rect 189 864 197 898
rect 147 739 197 864
rect 233 1411 241 1445
rect 275 1411 283 1445
rect 233 1034 283 1411
rect 233 1000 241 1034
rect 275 1000 283 1034
rect 233 966 283 1000
rect 233 932 241 966
rect 275 932 283 966
rect 233 898 283 932
rect 233 864 241 898
rect 275 864 283 898
rect 233 739 283 864
rect 319 1361 369 1445
rect 405 1411 413 1445
rect 447 1411 455 1445
rect 319 1327 327 1361
rect 361 1327 369 1361
rect 319 1034 369 1327
rect 319 1000 327 1034
rect 361 1000 369 1034
rect 319 966 369 1000
rect 319 932 327 966
rect 361 932 369 966
rect 319 898 369 932
rect 319 864 327 898
rect 361 864 369 898
rect 319 739 369 864
rect 233 605 283 689
rect 233 571 241 605
rect 275 571 283 605
rect 233 487 283 571
rect 233 185 283 269
rect 233 151 241 185
rect 275 151 283 185
rect 233 67 283 151
<< viali >>
rect 241 2839 275 2873
rect 241 2419 275 2453
rect 155 1663 189 1697
rect 241 1579 275 1613
rect 327 1663 361 1697
rect 413 1579 447 1613
rect 155 1327 189 1361
rect 241 1411 275 1445
rect 413 1411 447 1445
rect 327 1327 361 1361
rect 241 571 275 605
rect 241 151 275 185
<< metal1 >>
rect 138 2882 378 2884
rect 138 2830 146 2882
rect 198 2873 378 2882
rect 198 2839 241 2873
rect 275 2839 378 2873
rect 198 2830 378 2839
rect 138 2828 378 2830
rect 224 2462 464 2464
rect 224 2410 232 2462
rect 284 2410 464 2462
rect 224 2408 464 2410
rect 138 1706 378 1708
rect 138 1654 146 1706
rect 198 1697 378 1706
rect 198 1663 327 1697
rect 361 1663 378 1697
rect 198 1654 378 1663
rect 138 1652 378 1654
rect 224 1613 464 1624
rect 224 1579 241 1613
rect 275 1579 413 1613
rect 447 1579 464 1613
rect 224 1568 464 1579
rect 224 1445 464 1456
rect 224 1411 241 1445
rect 275 1411 413 1445
rect 447 1411 464 1445
rect 224 1400 464 1411
rect 138 1370 378 1372
rect 138 1318 146 1370
rect 198 1361 378 1370
rect 198 1327 327 1361
rect 361 1327 378 1361
rect 198 1318 378 1327
rect 138 1316 378 1318
rect 224 614 464 616
rect 224 562 232 614
rect 284 562 464 614
rect 224 560 464 562
rect 138 194 378 196
rect 138 142 146 194
rect 198 185 378 194
rect 198 151 241 185
rect 275 151 378 185
rect 198 142 378 151
rect 138 140 378 142
<< via1 >>
rect 146 2830 198 2882
rect 232 2453 284 2462
rect 232 2419 241 2453
rect 241 2419 275 2453
rect 275 2419 284 2453
rect 232 2410 284 2419
rect 146 1697 198 1706
rect 146 1663 155 1697
rect 155 1663 189 1697
rect 189 1663 198 1697
rect 146 1654 198 1663
rect 146 1361 198 1370
rect 146 1327 155 1361
rect 155 1327 189 1361
rect 189 1327 198 1361
rect 146 1318 198 1327
rect 232 605 284 614
rect 232 571 241 605
rect 241 571 275 605
rect 275 571 284 605
rect 232 562 284 571
rect 146 142 198 194
<< metal2 >>
rect 144 2882 200 2888
rect 144 2830 146 2882
rect 198 2830 200 2882
rect 144 1706 200 2830
rect 144 1654 146 1706
rect 198 1654 200 1706
rect 144 1648 200 1654
rect 230 2462 286 2468
rect 230 2410 232 2462
rect 284 2410 286 2462
rect 144 1370 200 1376
rect 144 1318 146 1370
rect 198 1318 200 1370
rect 144 194 200 1318
rect 230 614 286 2410
rect 230 562 232 614
rect 284 562 286 614
rect 230 556 286 562
rect 144 142 146 194
rect 198 142 200 194
rect 144 136 200 142
<< labels >>
flabel metal1 s 344 588 344 588 0 FreeSerif 0 0 0 0 A
flabel metal2 s 172 756 172 756 0 FreeSerif 0 0 0 0 VSS
flabel metal2 s 172 2268 172 2268 0 FreeSerif 0 0 0 0 VDD
flabel metal1 s 344 1428 344 1428 0 FreeSerif 0 0 0 0 Y
<< end >>
