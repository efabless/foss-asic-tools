magic
tech sky130A
magscale 1 2
timestamp 1622941822
<< nwell >>
rect -4940 40 4940 4500
<< pwell >>
rect -4940 -4500 4940 -40
<< mvpsubdiff >>
rect -4874 -118 4874 -106
rect -4874 -218 -4700 -118
rect 4700 -218 4874 -118
rect -4874 -230 4874 -218
rect -4874 -280 -4750 -230
rect -4874 -4260 -4862 -280
rect -4762 -4260 -4750 -280
rect -4874 -4310 -4750 -4260
rect 4750 -280 4874 -230
rect 4750 -4260 4762 -280
rect 4862 -4260 4874 -280
rect 4750 -4310 4874 -4260
rect -4874 -4322 4874 -4310
rect -4874 -4422 -4700 -4322
rect 4700 -4422 4874 -4322
rect -4874 -4434 4874 -4422
<< mvnsubdiff >>
rect -4874 4422 4874 4434
rect -4874 4322 -4700 4422
rect 4700 4322 4874 4422
rect -4874 4310 4874 4322
rect -4874 4260 -4750 4310
rect -4874 280 -4862 4260
rect -4762 280 -4750 4260
rect -4874 230 -4750 280
rect 4750 4260 4874 4310
rect 4750 280 4762 4260
rect 4862 280 4874 4260
rect 4750 230 4874 280
rect -4874 218 4874 230
rect -4874 118 -4700 218
rect 4700 118 4874 218
rect -4874 106 4874 118
<< mvpsubdiffcont >>
rect -4700 -218 4700 -118
rect -4862 -4260 -4762 -280
rect 4762 -4260 4862 -280
rect -4700 -4422 4700 -4322
<< mvnsubdiffcont >>
rect -4700 4322 4700 4422
rect -4862 280 -4762 4260
rect 4762 280 4862 4260
rect -4700 118 4700 218
<< locali >>
rect -4862 4260 -4762 4422
rect -4862 118 -4762 280
rect 4762 4260 4862 4422
rect 4762 118 4862 280
rect -4862 -280 -4762 -118
rect -4862 -4422 -4762 -4260
rect 4762 -280 4862 -118
rect 4762 -4422 4862 -4260
<< viali >>
rect -4762 4322 -4700 4422
rect -4700 4322 4700 4422
rect 4700 4322 4762 4422
rect -4862 423 -4762 4117
rect 4762 423 4862 4117
rect -4762 118 -4700 218
rect -4700 118 4700 218
rect 4700 118 4762 218
rect -4762 -218 -4700 -118
rect -4700 -218 4700 -118
rect 4700 -218 4762 -118
rect -4862 -4117 -4762 -423
rect 4762 -4117 4862 -423
rect -4762 -4422 -4700 -4322
rect -4700 -4422 4700 -4322
rect 4700 -4422 4762 -4322
<< metal1 >>
rect -4868 4422 4868 4428
rect -4868 4322 -4762 4422
rect 4762 4322 4868 4422
rect -4868 4316 4868 4322
rect -4868 4117 -4756 4316
rect -4868 423 -4862 4117
rect -4762 423 -4756 4117
rect -4156 4016 -4146 4316
rect 4146 4016 4156 4316
rect 4756 4117 4868 4316
rect -4868 224 -4756 423
rect 4756 423 4762 4117
rect 4862 423 4868 4117
rect 4756 224 4868 423
rect -4868 218 4868 224
rect -4868 118 -4762 218
rect 4762 118 4868 218
rect -4868 112 4868 118
rect -4868 -118 4868 -112
rect -4868 -218 -4762 -118
rect 4762 -218 4868 -118
rect -4868 -224 4868 -218
rect -4868 -423 -4756 -224
rect -4868 -4117 -4862 -423
rect -4762 -4117 -4756 -423
rect 4756 -423 4868 -224
rect -4868 -4316 -4756 -4117
rect -4156 -4316 -4146 -4016
rect 4146 -4316 4156 -4016
rect 4756 -4117 4762 -423
rect 4862 -4117 4868 -423
rect 4756 -4316 4868 -4117
rect -4868 -4322 4868 -4316
rect -4868 -4422 -4762 -4322
rect 4762 -4422 4868 -4322
rect -4868 -4428 4868 -4422
<< via1 >>
rect -4756 4016 -4156 4316
rect 4156 4016 4756 4316
rect -4756 -4316 -4156 -4016
rect 4156 -4316 4756 -4016
<< metal2 >>
rect -4756 4316 -4156 4326
rect -4756 4006 -4156 4016
rect 4156 4316 4756 4326
rect 4156 4006 4756 4016
rect -4756 -4016 -4156 -4006
rect -4756 -4326 -4156 -4316
rect 4156 -4016 4756 -4006
rect 4156 -4326 4756 -4316
<< via2 >>
rect -4756 4016 -4156 4316
rect 4156 4016 4756 4316
rect -4756 -4316 -4156 -4016
rect 4156 -4316 4756 -4016
<< metal3 >>
rect -4766 4316 -4146 4321
rect -4766 4016 -4756 4316
rect -4156 4016 -4146 4316
rect -4766 4011 -4146 4016
rect 4146 4316 4766 4321
rect 4146 4016 4156 4316
rect 4756 4016 4766 4316
rect 4146 4011 4766 4016
rect -4766 -4016 -4146 -4011
rect -4766 -4316 -4756 -4016
rect -4156 -4316 -4146 -4016
rect -4766 -4321 -4146 -4316
rect 4146 -4016 4766 -4011
rect 4146 -4316 4156 -4016
rect 4756 -4316 4766 -4016
rect 4146 -4321 4766 -4316
<< via3 >>
rect -4756 4016 -4156 4316
rect 4156 4016 4756 4316
rect -4756 -4316 -4156 -4016
rect 4156 -4316 4756 -4016
<< metal4 >>
rect -4940 4316 4940 4500
rect -4940 4016 -4756 4316
rect -4156 4016 4156 4316
rect 4756 4016 4940 4316
rect -4940 3700 4940 4016
rect -4940 -4016 4940 -3700
rect -4940 -4316 -4756 -4016
rect -4156 -4316 4156 -4016
rect 4756 -4316 4940 -4016
rect -4940 -4500 4940 -4316
use sky130_fd_pr__pfet_g5v0d10v5_8ATX2D  xm4
timestamp 1622941822
transform 1 0 0 0 1 3000
box -1514 -600 1514 600
use sky130_fd_pr__pfet_g5v0d10v5_ZD39PX  xm3
timestamp 1622941822
transform 1 0 0 0 1 1200
box -611 -600 611 600
use sky130_fd_pr__nfet_g5v0d10v5_7QEKRB  xm2
timestamp 1622941822
transform 1 0 0 0 1 -3000
box -2351 -588 2351 588
use sky130_fd_pr__nfet_g5v0d10v5_DQEKTK  xm1
timestamp 1622941822
transform 1 0 0 0 1 -1200
box -3899 -588 3899 588
<< labels >>
flabel metal4 -4940 3700 -4940 4500 3 FreeSans 480 0 0 0 vdd
port 1 e
flabel metal4 -4940 -4500 -4940 -3700 3 FreeSans 480 0 0 0 vss
port 2 e
<< properties >>
string FIXED_BBOX -4812 -4372 4812 -168
<< end >>
