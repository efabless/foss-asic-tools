magic
tech sky130A
magscale 1 2
timestamp 1678793193
<< nwell >>
rect 0 0 1204 2688
<< pwell >>
rect 1419 2382 2193 2658
rect 1325 1612 2287 1874
rect 1325 436 2287 698
<< nmos >>
rect 1404 1638 1434 1848
rect 1490 1638 1520 1848
rect 1576 1638 1606 1848
rect 1662 1638 1692 1848
rect 1748 1638 1778 1848
rect 1834 1638 1864 1848
rect 1920 1638 1950 1848
rect 2006 1638 2036 1848
rect 2092 1638 2122 1848
rect 2178 1638 2208 1848
rect 1404 462 1434 672
rect 1490 462 1520 672
rect 1576 462 1606 672
rect 1662 462 1692 672
rect 1748 462 1778 672
rect 1834 462 1864 672
rect 1920 462 1950 672
rect 2006 462 2036 672
rect 2092 462 2122 672
rect 2178 462 2208 672
<< pmos >>
rect 200 1659 230 1827
rect 286 1659 316 1827
rect 372 1659 402 1827
rect 458 1659 488 1827
rect 544 1659 574 1827
rect 630 1659 660 1827
rect 716 1659 746 1827
rect 802 1659 832 1827
rect 888 1659 918 1827
rect 974 1659 1004 1827
rect 200 483 230 651
rect 286 483 316 651
rect 372 483 402 651
rect 458 483 488 651
rect 544 483 574 651
rect 630 483 660 651
rect 716 483 746 651
rect 802 483 832 651
rect 888 483 918 651
rect 974 483 1004 651
<< ndiff >>
rect 1351 1824 1404 1848
rect 1351 1790 1359 1824
rect 1393 1790 1404 1824
rect 1351 1756 1404 1790
rect 1351 1722 1359 1756
rect 1393 1722 1404 1756
rect 1351 1688 1404 1722
rect 1351 1654 1359 1688
rect 1393 1654 1404 1688
rect 1351 1638 1404 1654
rect 1434 1824 1490 1848
rect 1434 1790 1445 1824
rect 1479 1790 1490 1824
rect 1434 1756 1490 1790
rect 1434 1722 1445 1756
rect 1479 1722 1490 1756
rect 1434 1688 1490 1722
rect 1434 1654 1445 1688
rect 1479 1654 1490 1688
rect 1434 1638 1490 1654
rect 1520 1824 1576 1848
rect 1520 1790 1531 1824
rect 1565 1790 1576 1824
rect 1520 1756 1576 1790
rect 1520 1722 1531 1756
rect 1565 1722 1576 1756
rect 1520 1688 1576 1722
rect 1520 1654 1531 1688
rect 1565 1654 1576 1688
rect 1520 1638 1576 1654
rect 1606 1824 1662 1848
rect 1606 1790 1617 1824
rect 1651 1790 1662 1824
rect 1606 1756 1662 1790
rect 1606 1722 1617 1756
rect 1651 1722 1662 1756
rect 1606 1688 1662 1722
rect 1606 1654 1617 1688
rect 1651 1654 1662 1688
rect 1606 1638 1662 1654
rect 1692 1824 1748 1848
rect 1692 1790 1703 1824
rect 1737 1790 1748 1824
rect 1692 1756 1748 1790
rect 1692 1722 1703 1756
rect 1737 1722 1748 1756
rect 1692 1688 1748 1722
rect 1692 1654 1703 1688
rect 1737 1654 1748 1688
rect 1692 1638 1748 1654
rect 1778 1824 1834 1848
rect 1778 1790 1789 1824
rect 1823 1790 1834 1824
rect 1778 1756 1834 1790
rect 1778 1722 1789 1756
rect 1823 1722 1834 1756
rect 1778 1688 1834 1722
rect 1778 1654 1789 1688
rect 1823 1654 1834 1688
rect 1778 1638 1834 1654
rect 1864 1824 1920 1848
rect 1864 1790 1875 1824
rect 1909 1790 1920 1824
rect 1864 1756 1920 1790
rect 1864 1722 1875 1756
rect 1909 1722 1920 1756
rect 1864 1688 1920 1722
rect 1864 1654 1875 1688
rect 1909 1654 1920 1688
rect 1864 1638 1920 1654
rect 1950 1824 2006 1848
rect 1950 1790 1961 1824
rect 1995 1790 2006 1824
rect 1950 1756 2006 1790
rect 1950 1722 1961 1756
rect 1995 1722 2006 1756
rect 1950 1688 2006 1722
rect 1950 1654 1961 1688
rect 1995 1654 2006 1688
rect 1950 1638 2006 1654
rect 2036 1824 2092 1848
rect 2036 1790 2047 1824
rect 2081 1790 2092 1824
rect 2036 1756 2092 1790
rect 2036 1722 2047 1756
rect 2081 1722 2092 1756
rect 2036 1688 2092 1722
rect 2036 1654 2047 1688
rect 2081 1654 2092 1688
rect 2036 1638 2092 1654
rect 2122 1824 2178 1848
rect 2122 1790 2133 1824
rect 2167 1790 2178 1824
rect 2122 1756 2178 1790
rect 2122 1722 2133 1756
rect 2167 1722 2178 1756
rect 2122 1688 2178 1722
rect 2122 1654 2133 1688
rect 2167 1654 2178 1688
rect 2122 1638 2178 1654
rect 2208 1824 2261 1848
rect 2208 1790 2219 1824
rect 2253 1790 2261 1824
rect 2208 1756 2261 1790
rect 2208 1722 2219 1756
rect 2253 1722 2261 1756
rect 2208 1688 2261 1722
rect 2208 1654 2219 1688
rect 2253 1654 2261 1688
rect 2208 1638 2261 1654
rect 1351 648 1404 672
rect 1351 614 1359 648
rect 1393 614 1404 648
rect 1351 580 1404 614
rect 1351 546 1359 580
rect 1393 546 1404 580
rect 1351 512 1404 546
rect 1351 478 1359 512
rect 1393 478 1404 512
rect 1351 462 1404 478
rect 1434 648 1490 672
rect 1434 614 1445 648
rect 1479 614 1490 648
rect 1434 580 1490 614
rect 1434 546 1445 580
rect 1479 546 1490 580
rect 1434 512 1490 546
rect 1434 478 1445 512
rect 1479 478 1490 512
rect 1434 462 1490 478
rect 1520 648 1576 672
rect 1520 614 1531 648
rect 1565 614 1576 648
rect 1520 580 1576 614
rect 1520 546 1531 580
rect 1565 546 1576 580
rect 1520 512 1576 546
rect 1520 478 1531 512
rect 1565 478 1576 512
rect 1520 462 1576 478
rect 1606 648 1662 672
rect 1606 614 1617 648
rect 1651 614 1662 648
rect 1606 580 1662 614
rect 1606 546 1617 580
rect 1651 546 1662 580
rect 1606 512 1662 546
rect 1606 478 1617 512
rect 1651 478 1662 512
rect 1606 462 1662 478
rect 1692 648 1748 672
rect 1692 614 1703 648
rect 1737 614 1748 648
rect 1692 580 1748 614
rect 1692 546 1703 580
rect 1737 546 1748 580
rect 1692 512 1748 546
rect 1692 478 1703 512
rect 1737 478 1748 512
rect 1692 462 1748 478
rect 1778 648 1834 672
rect 1778 614 1789 648
rect 1823 614 1834 648
rect 1778 580 1834 614
rect 1778 546 1789 580
rect 1823 546 1834 580
rect 1778 512 1834 546
rect 1778 478 1789 512
rect 1823 478 1834 512
rect 1778 462 1834 478
rect 1864 648 1920 672
rect 1864 614 1875 648
rect 1909 614 1920 648
rect 1864 580 1920 614
rect 1864 546 1875 580
rect 1909 546 1920 580
rect 1864 512 1920 546
rect 1864 478 1875 512
rect 1909 478 1920 512
rect 1864 462 1920 478
rect 1950 648 2006 672
rect 1950 614 1961 648
rect 1995 614 2006 648
rect 1950 580 2006 614
rect 1950 546 1961 580
rect 1995 546 2006 580
rect 1950 512 2006 546
rect 1950 478 1961 512
rect 1995 478 2006 512
rect 1950 462 2006 478
rect 2036 648 2092 672
rect 2036 614 2047 648
rect 2081 614 2092 648
rect 2036 580 2092 614
rect 2036 546 2047 580
rect 2081 546 2092 580
rect 2036 512 2092 546
rect 2036 478 2047 512
rect 2081 478 2092 512
rect 2036 462 2092 478
rect 2122 648 2178 672
rect 2122 614 2133 648
rect 2167 614 2178 648
rect 2122 580 2178 614
rect 2122 546 2133 580
rect 2167 546 2178 580
rect 2122 512 2178 546
rect 2122 478 2133 512
rect 2167 478 2178 512
rect 2122 462 2178 478
rect 2208 648 2261 672
rect 2208 614 2219 648
rect 2253 614 2261 648
rect 2208 580 2261 614
rect 2208 546 2219 580
rect 2253 546 2261 580
rect 2208 512 2261 546
rect 2208 478 2219 512
rect 2253 478 2261 512
rect 2208 462 2261 478
<< pdiff >>
rect 147 1777 200 1827
rect 147 1743 155 1777
rect 189 1743 200 1777
rect 147 1709 200 1743
rect 147 1675 155 1709
rect 189 1675 200 1709
rect 147 1659 200 1675
rect 230 1777 286 1827
rect 230 1743 241 1777
rect 275 1743 286 1777
rect 230 1709 286 1743
rect 230 1675 241 1709
rect 275 1675 286 1709
rect 230 1659 286 1675
rect 316 1777 372 1827
rect 316 1743 327 1777
rect 361 1743 372 1777
rect 316 1709 372 1743
rect 316 1675 327 1709
rect 361 1675 372 1709
rect 316 1659 372 1675
rect 402 1777 458 1827
rect 402 1743 413 1777
rect 447 1743 458 1777
rect 402 1709 458 1743
rect 402 1675 413 1709
rect 447 1675 458 1709
rect 402 1659 458 1675
rect 488 1777 544 1827
rect 488 1743 499 1777
rect 533 1743 544 1777
rect 488 1709 544 1743
rect 488 1675 499 1709
rect 533 1675 544 1709
rect 488 1659 544 1675
rect 574 1777 630 1827
rect 574 1743 585 1777
rect 619 1743 630 1777
rect 574 1709 630 1743
rect 574 1675 585 1709
rect 619 1675 630 1709
rect 574 1659 630 1675
rect 660 1777 716 1827
rect 660 1743 671 1777
rect 705 1743 716 1777
rect 660 1709 716 1743
rect 660 1675 671 1709
rect 705 1675 716 1709
rect 660 1659 716 1675
rect 746 1777 802 1827
rect 746 1743 757 1777
rect 791 1743 802 1777
rect 746 1709 802 1743
rect 746 1675 757 1709
rect 791 1675 802 1709
rect 746 1659 802 1675
rect 832 1777 888 1827
rect 832 1743 843 1777
rect 877 1743 888 1777
rect 832 1709 888 1743
rect 832 1675 843 1709
rect 877 1675 888 1709
rect 832 1659 888 1675
rect 918 1777 974 1827
rect 918 1743 929 1777
rect 963 1743 974 1777
rect 918 1709 974 1743
rect 918 1675 929 1709
rect 963 1675 974 1709
rect 918 1659 974 1675
rect 1004 1777 1057 1827
rect 1004 1743 1015 1777
rect 1049 1743 1057 1777
rect 1004 1709 1057 1743
rect 1004 1675 1015 1709
rect 1049 1675 1057 1709
rect 1004 1659 1057 1675
rect 147 601 200 651
rect 147 567 155 601
rect 189 567 200 601
rect 147 533 200 567
rect 147 499 155 533
rect 189 499 200 533
rect 147 483 200 499
rect 230 601 286 651
rect 230 567 241 601
rect 275 567 286 601
rect 230 533 286 567
rect 230 499 241 533
rect 275 499 286 533
rect 230 483 286 499
rect 316 601 372 651
rect 316 567 327 601
rect 361 567 372 601
rect 316 533 372 567
rect 316 499 327 533
rect 361 499 372 533
rect 316 483 372 499
rect 402 601 458 651
rect 402 567 413 601
rect 447 567 458 601
rect 402 533 458 567
rect 402 499 413 533
rect 447 499 458 533
rect 402 483 458 499
rect 488 601 544 651
rect 488 567 499 601
rect 533 567 544 601
rect 488 533 544 567
rect 488 499 499 533
rect 533 499 544 533
rect 488 483 544 499
rect 574 601 630 651
rect 574 567 585 601
rect 619 567 630 601
rect 574 533 630 567
rect 574 499 585 533
rect 619 499 630 533
rect 574 483 630 499
rect 660 601 716 651
rect 660 567 671 601
rect 705 567 716 601
rect 660 533 716 567
rect 660 499 671 533
rect 705 499 716 533
rect 660 483 716 499
rect 746 601 802 651
rect 746 567 757 601
rect 791 567 802 601
rect 746 533 802 567
rect 746 499 757 533
rect 791 499 802 533
rect 746 483 802 499
rect 832 601 888 651
rect 832 567 843 601
rect 877 567 888 601
rect 832 533 888 567
rect 832 499 843 533
rect 877 499 888 533
rect 832 483 888 499
rect 918 601 974 651
rect 918 567 929 601
rect 963 567 974 601
rect 918 533 974 567
rect 918 499 929 533
rect 963 499 974 533
rect 918 483 974 499
rect 1004 601 1057 651
rect 1004 567 1015 601
rect 1049 567 1057 601
rect 1004 533 1057 567
rect 1004 499 1015 533
rect 1049 499 1057 533
rect 1004 483 1057 499
<< ndiffc >>
rect 1359 1790 1393 1824
rect 1359 1722 1393 1756
rect 1359 1654 1393 1688
rect 1445 1790 1479 1824
rect 1445 1722 1479 1756
rect 1445 1654 1479 1688
rect 1531 1790 1565 1824
rect 1531 1722 1565 1756
rect 1531 1654 1565 1688
rect 1617 1790 1651 1824
rect 1617 1722 1651 1756
rect 1617 1654 1651 1688
rect 1703 1790 1737 1824
rect 1703 1722 1737 1756
rect 1703 1654 1737 1688
rect 1789 1790 1823 1824
rect 1789 1722 1823 1756
rect 1789 1654 1823 1688
rect 1875 1790 1909 1824
rect 1875 1722 1909 1756
rect 1875 1654 1909 1688
rect 1961 1790 1995 1824
rect 1961 1722 1995 1756
rect 1961 1654 1995 1688
rect 2047 1790 2081 1824
rect 2047 1722 2081 1756
rect 2047 1654 2081 1688
rect 2133 1790 2167 1824
rect 2133 1722 2167 1756
rect 2133 1654 2167 1688
rect 2219 1790 2253 1824
rect 2219 1722 2253 1756
rect 2219 1654 2253 1688
rect 1359 614 1393 648
rect 1359 546 1393 580
rect 1359 478 1393 512
rect 1445 614 1479 648
rect 1445 546 1479 580
rect 1445 478 1479 512
rect 1531 614 1565 648
rect 1531 546 1565 580
rect 1531 478 1565 512
rect 1617 614 1651 648
rect 1617 546 1651 580
rect 1617 478 1651 512
rect 1703 614 1737 648
rect 1703 546 1737 580
rect 1703 478 1737 512
rect 1789 614 1823 648
rect 1789 546 1823 580
rect 1789 478 1823 512
rect 1875 614 1909 648
rect 1875 546 1909 580
rect 1875 478 1909 512
rect 1961 614 1995 648
rect 1961 546 1995 580
rect 1961 478 1995 512
rect 2047 614 2081 648
rect 2047 546 2081 580
rect 2047 478 2081 512
rect 2133 614 2167 648
rect 2133 546 2167 580
rect 2133 478 2167 512
rect 2219 614 2253 648
rect 2219 546 2253 580
rect 2219 478 2253 512
<< pdiffc >>
rect 155 1743 189 1777
rect 155 1675 189 1709
rect 241 1743 275 1777
rect 241 1675 275 1709
rect 327 1743 361 1777
rect 327 1675 361 1709
rect 413 1743 447 1777
rect 413 1675 447 1709
rect 499 1743 533 1777
rect 499 1675 533 1709
rect 585 1743 619 1777
rect 585 1675 619 1709
rect 671 1743 705 1777
rect 671 1675 705 1709
rect 757 1743 791 1777
rect 757 1675 791 1709
rect 843 1743 877 1777
rect 843 1675 877 1709
rect 929 1743 963 1777
rect 929 1675 963 1709
rect 1015 1743 1049 1777
rect 1015 1675 1049 1709
rect 155 567 189 601
rect 155 499 189 533
rect 241 567 275 601
rect 241 499 275 533
rect 327 567 361 601
rect 327 499 361 533
rect 413 567 447 601
rect 413 499 447 533
rect 499 567 533 601
rect 499 499 533 533
rect 585 567 619 601
rect 585 499 619 533
rect 671 567 705 601
rect 671 499 705 533
rect 757 567 791 601
rect 757 499 791 533
rect 843 567 877 601
rect 843 499 877 533
rect 929 567 963 601
rect 929 499 963 533
rect 1015 567 1049 601
rect 1015 499 1049 533
<< psubdiff >>
rect 1445 2537 1479 2632
rect 1445 2408 1479 2503
rect 1617 2537 1651 2632
rect 1617 2408 1651 2503
rect 1789 2537 1823 2632
rect 1789 2408 1823 2503
rect 1961 2537 1995 2632
rect 1961 2408 1995 2503
rect 2133 2537 2167 2632
rect 2133 2408 2167 2503
<< nsubdiff >>
rect 241 2537 275 2632
rect 241 2408 275 2503
rect 413 2537 447 2632
rect 413 2408 447 2503
rect 585 2537 619 2632
rect 585 2408 619 2503
rect 757 2537 791 2632
rect 757 2408 791 2503
rect 929 2537 963 2632
rect 929 2408 963 2503
<< psubdiffcont >>
rect 1445 2503 1479 2537
rect 1617 2503 1651 2537
rect 1789 2503 1823 2537
rect 1961 2503 1995 2537
rect 2133 2503 2167 2537
<< nsubdiffcont >>
rect 241 2503 275 2537
rect 413 2503 447 2537
rect 585 2503 619 2537
rect 757 2503 791 2537
rect 929 2503 963 2537
<< poly >>
rect 200 2117 316 2127
rect 200 2083 241 2117
rect 275 2083 316 2117
rect 200 2073 316 2083
rect 200 1827 230 2073
rect 286 1827 316 2073
rect 372 2117 488 2127
rect 372 2083 413 2117
rect 447 2083 488 2117
rect 372 2073 488 2083
rect 372 1827 402 2073
rect 458 1827 488 2073
rect 544 2117 660 2127
rect 544 2083 585 2117
rect 619 2083 660 2117
rect 544 2073 660 2083
rect 544 1827 574 2073
rect 630 1827 660 2073
rect 716 2117 832 2127
rect 716 2083 757 2117
rect 791 2083 832 2117
rect 716 2073 832 2083
rect 716 1827 746 2073
rect 802 1827 832 2073
rect 888 2117 1004 2127
rect 888 2083 929 2117
rect 963 2083 1004 2117
rect 888 2073 1004 2083
rect 888 1827 918 2073
rect 974 1827 1004 2073
rect 1404 2117 1520 2127
rect 1404 2083 1445 2117
rect 1479 2083 1520 2117
rect 1404 2073 1520 2083
rect 1404 1848 1434 2073
rect 1490 1848 1520 2073
rect 1576 2117 1692 2127
rect 1576 2083 1617 2117
rect 1651 2083 1692 2117
rect 1576 2073 1692 2083
rect 1576 1848 1606 2073
rect 1662 1848 1692 2073
rect 1748 2117 1864 2127
rect 1748 2083 1789 2117
rect 1823 2083 1864 2117
rect 1748 2073 1864 2083
rect 1748 1848 1778 2073
rect 1834 1848 1864 2073
rect 1920 2117 2036 2127
rect 1920 2083 1961 2117
rect 1995 2083 2036 2117
rect 1920 2073 2036 2083
rect 1920 1848 1950 2073
rect 2006 1848 2036 2073
rect 2092 2117 2208 2127
rect 2092 2083 2133 2117
rect 2167 2083 2208 2117
rect 2092 2073 2208 2083
rect 2092 1848 2122 2073
rect 2178 1848 2208 2073
rect 200 1428 230 1659
rect 286 1428 316 1659
rect 372 1428 402 1659
rect 458 1428 488 1659
rect 544 1428 574 1659
rect 630 1428 660 1659
rect 716 1428 746 1659
rect 802 1428 832 1659
rect 888 1428 918 1659
rect 974 1428 1004 1659
rect 1404 1428 1434 1638
rect 1490 1428 1520 1638
rect 1576 1428 1606 1638
rect 1662 1428 1692 1638
rect 1748 1428 1778 1638
rect 1834 1428 1864 1638
rect 1920 1428 1950 1638
rect 2006 1428 2036 1638
rect 2092 1428 2122 1638
rect 2178 1428 2208 1638
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 651 230 897
rect 286 651 316 897
rect 372 941 488 951
rect 372 907 413 941
rect 447 907 488 941
rect 372 897 488 907
rect 372 651 402 897
rect 458 651 488 897
rect 544 941 660 951
rect 544 907 585 941
rect 619 907 660 941
rect 544 897 660 907
rect 544 651 574 897
rect 630 651 660 897
rect 716 941 832 951
rect 716 907 757 941
rect 791 907 832 941
rect 716 897 832 907
rect 716 651 746 897
rect 802 651 832 897
rect 888 941 1004 951
rect 888 907 929 941
rect 963 907 1004 941
rect 888 897 1004 907
rect 888 651 918 897
rect 974 651 1004 897
rect 1404 941 1520 951
rect 1404 907 1445 941
rect 1479 907 1520 941
rect 1404 897 1520 907
rect 1404 672 1434 897
rect 1490 672 1520 897
rect 1576 941 1692 951
rect 1576 907 1617 941
rect 1651 907 1692 941
rect 1576 897 1692 907
rect 1576 672 1606 897
rect 1662 672 1692 897
rect 1748 941 1864 951
rect 1748 907 1789 941
rect 1823 907 1864 941
rect 1748 897 1864 907
rect 1748 672 1778 897
rect 1834 672 1864 897
rect 1920 941 2036 951
rect 1920 907 1961 941
rect 1995 907 2036 941
rect 1920 897 2036 907
rect 1920 672 1950 897
rect 2006 672 2036 897
rect 2092 941 2208 951
rect 2092 907 2133 941
rect 2167 907 2208 941
rect 2092 897 2208 907
rect 2092 672 2122 897
rect 2178 672 2208 897
rect 200 252 230 483
rect 286 252 316 483
rect 372 252 402 483
rect 458 252 488 483
rect 544 252 574 483
rect 630 252 660 483
rect 716 252 746 483
rect 802 252 832 483
rect 888 252 918 483
rect 974 252 1004 483
rect 1404 252 1434 462
rect 1490 252 1520 462
rect 1576 252 1606 462
rect 1662 252 1692 462
rect 1748 252 1778 462
rect 1834 252 1864 462
rect 1920 252 1950 462
rect 2006 252 2036 462
rect 2092 252 2122 462
rect 2178 252 2208 462
<< polycont >>
rect 241 2083 275 2117
rect 413 2083 447 2117
rect 585 2083 619 2117
rect 757 2083 791 2117
rect 929 2083 963 2117
rect 1445 2083 1479 2117
rect 1617 2083 1651 2117
rect 1789 2083 1823 2117
rect 1961 2083 1995 2117
rect 2133 2083 2167 2117
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
rect 1445 907 1479 941
rect 1617 907 1651 941
rect 1789 907 1823 941
rect 1961 907 1995 941
rect 2133 907 2167 941
<< locali >>
rect 233 2537 283 2621
rect 233 2503 241 2537
rect 275 2503 283 2537
rect 233 2419 283 2503
rect 405 2537 455 2621
rect 405 2503 413 2537
rect 447 2503 455 2537
rect 405 2419 455 2503
rect 577 2537 627 2621
rect 577 2503 585 2537
rect 619 2503 627 2537
rect 577 2419 627 2503
rect 749 2537 799 2621
rect 749 2503 757 2537
rect 791 2503 799 2537
rect 749 2419 799 2503
rect 921 2537 971 2621
rect 921 2503 929 2537
rect 963 2503 971 2537
rect 921 2419 971 2503
rect 1437 2537 1487 2621
rect 1437 2503 1445 2537
rect 1479 2503 1487 2537
rect 1437 2419 1487 2503
rect 1609 2537 1659 2621
rect 1609 2503 1617 2537
rect 1651 2503 1659 2537
rect 1609 2419 1659 2503
rect 1781 2537 1831 2621
rect 1781 2503 1789 2537
rect 1823 2503 1831 2537
rect 1781 2419 1831 2503
rect 1953 2537 2003 2621
rect 1953 2503 1961 2537
rect 1995 2503 2003 2537
rect 1953 2419 2003 2503
rect 2125 2537 2175 2621
rect 2125 2503 2133 2537
rect 2167 2503 2175 2537
rect 2125 2419 2175 2503
rect 233 2117 283 2201
rect 233 2083 241 2117
rect 275 2083 283 2117
rect 233 1999 283 2083
rect 405 2117 455 2201
rect 405 2083 413 2117
rect 447 2083 455 2117
rect 405 1999 455 2083
rect 577 2117 627 2201
rect 577 2083 585 2117
rect 619 2083 627 2117
rect 577 1999 627 2083
rect 749 2117 799 2201
rect 749 2083 757 2117
rect 791 2083 799 2117
rect 749 1999 799 2083
rect 921 2117 971 2201
rect 921 2083 929 2117
rect 963 2083 971 2117
rect 921 1999 971 2083
rect 1437 2117 1487 2201
rect 1437 2083 1445 2117
rect 1479 2083 1487 2117
rect 1437 1999 1487 2083
rect 1609 2117 1659 2201
rect 1609 2083 1617 2117
rect 1651 2083 1659 2117
rect 1609 1999 1659 2083
rect 1781 2117 1831 2201
rect 1781 2083 1789 2117
rect 1823 2083 1831 2117
rect 1781 1999 1831 2083
rect 1953 2117 2003 2201
rect 1953 2083 1961 2117
rect 1995 2083 2003 2117
rect 1953 1999 2003 2083
rect 2125 2117 2175 2201
rect 2125 2083 2133 2117
rect 2167 2083 2175 2117
rect 2125 1999 2175 2083
rect 147 1777 197 1949
rect 147 1743 155 1777
rect 189 1743 197 1777
rect 147 1709 197 1743
rect 147 1675 155 1709
rect 189 1675 197 1709
rect 147 1361 197 1675
rect 147 1327 155 1361
rect 189 1327 197 1361
rect 147 1243 197 1327
rect 233 1777 283 1949
rect 233 1743 241 1777
rect 275 1743 283 1777
rect 233 1709 283 1743
rect 233 1675 241 1709
rect 275 1675 283 1709
rect 233 1277 283 1675
rect 233 1243 241 1277
rect 275 1243 283 1277
rect 319 1777 369 1949
rect 319 1743 327 1777
rect 361 1743 369 1777
rect 319 1709 369 1743
rect 319 1675 327 1709
rect 361 1675 369 1709
rect 319 1361 369 1675
rect 319 1327 327 1361
rect 361 1327 369 1361
rect 319 1243 369 1327
rect 405 1777 455 1949
rect 405 1743 413 1777
rect 447 1743 455 1777
rect 405 1709 455 1743
rect 405 1675 413 1709
rect 447 1675 455 1709
rect 405 1277 455 1675
rect 405 1243 413 1277
rect 447 1243 455 1277
rect 491 1777 541 1949
rect 491 1743 499 1777
rect 533 1743 541 1777
rect 491 1709 541 1743
rect 491 1675 499 1709
rect 533 1675 541 1709
rect 491 1361 541 1675
rect 491 1327 499 1361
rect 533 1327 541 1361
rect 491 1243 541 1327
rect 577 1777 627 1949
rect 577 1743 585 1777
rect 619 1743 627 1777
rect 577 1709 627 1743
rect 577 1675 585 1709
rect 619 1675 627 1709
rect 577 1277 627 1675
rect 577 1243 585 1277
rect 619 1243 627 1277
rect 663 1777 713 1949
rect 663 1743 671 1777
rect 705 1743 713 1777
rect 663 1709 713 1743
rect 663 1675 671 1709
rect 705 1675 713 1709
rect 663 1361 713 1675
rect 663 1327 671 1361
rect 705 1327 713 1361
rect 663 1243 713 1327
rect 749 1777 799 1949
rect 749 1743 757 1777
rect 791 1743 799 1777
rect 749 1709 799 1743
rect 749 1675 757 1709
rect 791 1675 799 1709
rect 749 1277 799 1675
rect 749 1243 757 1277
rect 791 1243 799 1277
rect 835 1777 885 1949
rect 835 1743 843 1777
rect 877 1743 885 1777
rect 835 1709 885 1743
rect 835 1675 843 1709
rect 877 1675 885 1709
rect 835 1361 885 1675
rect 835 1327 843 1361
rect 877 1327 885 1361
rect 835 1243 885 1327
rect 921 1777 971 1949
rect 921 1743 929 1777
rect 963 1743 971 1777
rect 921 1709 971 1743
rect 921 1675 929 1709
rect 963 1675 971 1709
rect 921 1277 971 1675
rect 921 1243 929 1277
rect 963 1243 971 1277
rect 1007 1777 1057 1949
rect 1007 1743 1015 1777
rect 1049 1743 1057 1777
rect 1007 1709 1057 1743
rect 1007 1675 1015 1709
rect 1049 1675 1057 1709
rect 1007 1361 1057 1675
rect 1007 1327 1015 1361
rect 1049 1327 1057 1361
rect 1007 1243 1057 1327
rect 1351 1824 1401 1949
rect 1351 1790 1359 1824
rect 1393 1790 1401 1824
rect 1351 1756 1401 1790
rect 1351 1722 1359 1756
rect 1393 1722 1401 1756
rect 1351 1688 1401 1722
rect 1351 1654 1359 1688
rect 1393 1654 1401 1688
rect 1351 1361 1401 1654
rect 1351 1327 1359 1361
rect 1393 1327 1401 1361
rect 1351 1243 1401 1327
rect 1437 1824 1487 1949
rect 1437 1790 1445 1824
rect 1479 1790 1487 1824
rect 1437 1756 1487 1790
rect 1437 1722 1445 1756
rect 1479 1722 1487 1756
rect 1437 1688 1487 1722
rect 1437 1654 1445 1688
rect 1479 1654 1487 1688
rect 1437 1277 1487 1654
rect 1437 1243 1445 1277
rect 1479 1243 1487 1277
rect 1523 1824 1573 1949
rect 1523 1790 1531 1824
rect 1565 1790 1573 1824
rect 1523 1756 1573 1790
rect 1523 1722 1531 1756
rect 1565 1722 1573 1756
rect 1523 1688 1573 1722
rect 1523 1654 1531 1688
rect 1565 1654 1573 1688
rect 1523 1361 1573 1654
rect 1523 1327 1531 1361
rect 1565 1327 1573 1361
rect 1523 1243 1573 1327
rect 1609 1824 1659 1949
rect 1609 1790 1617 1824
rect 1651 1790 1659 1824
rect 1609 1756 1659 1790
rect 1609 1722 1617 1756
rect 1651 1722 1659 1756
rect 1609 1688 1659 1722
rect 1609 1654 1617 1688
rect 1651 1654 1659 1688
rect 1609 1277 1659 1654
rect 1609 1243 1617 1277
rect 1651 1243 1659 1277
rect 1695 1824 1745 1949
rect 1695 1790 1703 1824
rect 1737 1790 1745 1824
rect 1695 1756 1745 1790
rect 1695 1722 1703 1756
rect 1737 1722 1745 1756
rect 1695 1688 1745 1722
rect 1695 1654 1703 1688
rect 1737 1654 1745 1688
rect 1695 1361 1745 1654
rect 1695 1327 1703 1361
rect 1737 1327 1745 1361
rect 1695 1243 1745 1327
rect 1781 1824 1831 1949
rect 1781 1790 1789 1824
rect 1823 1790 1831 1824
rect 1781 1756 1831 1790
rect 1781 1722 1789 1756
rect 1823 1722 1831 1756
rect 1781 1688 1831 1722
rect 1781 1654 1789 1688
rect 1823 1654 1831 1688
rect 1781 1277 1831 1654
rect 1781 1243 1789 1277
rect 1823 1243 1831 1277
rect 1867 1824 1917 1949
rect 1867 1790 1875 1824
rect 1909 1790 1917 1824
rect 1867 1756 1917 1790
rect 1867 1722 1875 1756
rect 1909 1722 1917 1756
rect 1867 1688 1917 1722
rect 1867 1654 1875 1688
rect 1909 1654 1917 1688
rect 1867 1361 1917 1654
rect 1867 1327 1875 1361
rect 1909 1327 1917 1361
rect 1867 1243 1917 1327
rect 1953 1824 2003 1949
rect 1953 1790 1961 1824
rect 1995 1790 2003 1824
rect 1953 1756 2003 1790
rect 1953 1722 1961 1756
rect 1995 1722 2003 1756
rect 1953 1688 2003 1722
rect 1953 1654 1961 1688
rect 1995 1654 2003 1688
rect 1953 1277 2003 1654
rect 1953 1243 1961 1277
rect 1995 1243 2003 1277
rect 2039 1824 2089 1949
rect 2039 1790 2047 1824
rect 2081 1790 2089 1824
rect 2039 1756 2089 1790
rect 2039 1722 2047 1756
rect 2081 1722 2089 1756
rect 2039 1688 2089 1722
rect 2039 1654 2047 1688
rect 2081 1654 2089 1688
rect 2039 1361 2089 1654
rect 2039 1327 2047 1361
rect 2081 1327 2089 1361
rect 2039 1243 2089 1327
rect 2125 1824 2175 1949
rect 2125 1790 2133 1824
rect 2167 1790 2175 1824
rect 2125 1756 2175 1790
rect 2125 1722 2133 1756
rect 2167 1722 2175 1756
rect 2125 1688 2175 1722
rect 2125 1654 2133 1688
rect 2167 1654 2175 1688
rect 2125 1277 2175 1654
rect 2125 1243 2133 1277
rect 2167 1243 2175 1277
rect 2211 1824 2261 1949
rect 2211 1790 2219 1824
rect 2253 1790 2261 1824
rect 2211 1756 2261 1790
rect 2211 1722 2219 1756
rect 2253 1722 2261 1756
rect 2211 1688 2261 1722
rect 2211 1654 2219 1688
rect 2253 1654 2261 1688
rect 2211 1361 2261 1654
rect 2211 1327 2219 1361
rect 2253 1327 2261 1361
rect 2211 1243 2261 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 405 941 455 1025
rect 405 907 413 941
rect 447 907 455 941
rect 405 823 455 907
rect 577 941 627 1025
rect 577 907 585 941
rect 619 907 627 941
rect 577 823 627 907
rect 749 941 799 1025
rect 749 907 757 941
rect 791 907 799 941
rect 749 823 799 907
rect 921 941 971 1025
rect 921 907 929 941
rect 963 907 971 941
rect 921 823 971 907
rect 1437 941 1487 1025
rect 1437 907 1445 941
rect 1479 907 1487 941
rect 1437 823 1487 907
rect 1609 941 1659 1025
rect 1609 907 1617 941
rect 1651 907 1659 941
rect 1609 823 1659 907
rect 1781 941 1831 1025
rect 1781 907 1789 941
rect 1823 907 1831 941
rect 1781 823 1831 907
rect 1953 941 2003 1025
rect 1953 907 1961 941
rect 1995 907 2003 941
rect 1953 823 2003 907
rect 2125 941 2175 1025
rect 2125 907 2133 941
rect 2167 907 2175 941
rect 2125 823 2175 907
rect 147 601 197 773
rect 147 567 155 601
rect 189 567 197 601
rect 147 533 197 567
rect 147 499 155 533
rect 189 499 197 533
rect 147 185 197 499
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 601 283 773
rect 233 567 241 601
rect 275 567 283 601
rect 233 533 283 567
rect 233 499 241 533
rect 275 499 283 533
rect 233 101 283 499
rect 233 67 241 101
rect 275 67 283 101
rect 319 601 369 773
rect 319 567 327 601
rect 361 567 369 601
rect 319 533 369 567
rect 319 499 327 533
rect 361 499 369 533
rect 319 185 369 499
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
rect 405 601 455 773
rect 405 567 413 601
rect 447 567 455 601
rect 405 533 455 567
rect 405 499 413 533
rect 447 499 455 533
rect 405 101 455 499
rect 405 67 413 101
rect 447 67 455 101
rect 491 601 541 773
rect 491 567 499 601
rect 533 567 541 601
rect 491 533 541 567
rect 491 499 499 533
rect 533 499 541 533
rect 491 185 541 499
rect 491 151 499 185
rect 533 151 541 185
rect 491 67 541 151
rect 577 601 627 773
rect 577 567 585 601
rect 619 567 627 601
rect 577 533 627 567
rect 577 499 585 533
rect 619 499 627 533
rect 577 101 627 499
rect 577 67 585 101
rect 619 67 627 101
rect 663 601 713 773
rect 663 567 671 601
rect 705 567 713 601
rect 663 533 713 567
rect 663 499 671 533
rect 705 499 713 533
rect 663 185 713 499
rect 663 151 671 185
rect 705 151 713 185
rect 663 67 713 151
rect 749 601 799 773
rect 749 567 757 601
rect 791 567 799 601
rect 749 533 799 567
rect 749 499 757 533
rect 791 499 799 533
rect 749 101 799 499
rect 749 67 757 101
rect 791 67 799 101
rect 835 601 885 773
rect 835 567 843 601
rect 877 567 885 601
rect 835 533 885 567
rect 835 499 843 533
rect 877 499 885 533
rect 835 185 885 499
rect 835 151 843 185
rect 877 151 885 185
rect 835 67 885 151
rect 921 601 971 773
rect 921 567 929 601
rect 963 567 971 601
rect 921 533 971 567
rect 921 499 929 533
rect 963 499 971 533
rect 921 101 971 499
rect 921 67 929 101
rect 963 67 971 101
rect 1007 601 1057 773
rect 1007 567 1015 601
rect 1049 567 1057 601
rect 1007 533 1057 567
rect 1007 499 1015 533
rect 1049 499 1057 533
rect 1007 185 1057 499
rect 1007 151 1015 185
rect 1049 151 1057 185
rect 1007 67 1057 151
rect 1351 648 1401 773
rect 1351 614 1359 648
rect 1393 614 1401 648
rect 1351 580 1401 614
rect 1351 546 1359 580
rect 1393 546 1401 580
rect 1351 512 1401 546
rect 1351 478 1359 512
rect 1393 478 1401 512
rect 1351 185 1401 478
rect 1351 151 1359 185
rect 1393 151 1401 185
rect 1351 67 1401 151
rect 1437 648 1487 773
rect 1437 614 1445 648
rect 1479 614 1487 648
rect 1437 580 1487 614
rect 1437 546 1445 580
rect 1479 546 1487 580
rect 1437 512 1487 546
rect 1437 478 1445 512
rect 1479 478 1487 512
rect 1437 101 1487 478
rect 1437 67 1445 101
rect 1479 67 1487 101
rect 1523 648 1573 773
rect 1523 614 1531 648
rect 1565 614 1573 648
rect 1523 580 1573 614
rect 1523 546 1531 580
rect 1565 546 1573 580
rect 1523 512 1573 546
rect 1523 478 1531 512
rect 1565 478 1573 512
rect 1523 185 1573 478
rect 1523 151 1531 185
rect 1565 151 1573 185
rect 1523 67 1573 151
rect 1609 648 1659 773
rect 1609 614 1617 648
rect 1651 614 1659 648
rect 1609 580 1659 614
rect 1609 546 1617 580
rect 1651 546 1659 580
rect 1609 512 1659 546
rect 1609 478 1617 512
rect 1651 478 1659 512
rect 1609 101 1659 478
rect 1609 67 1617 101
rect 1651 67 1659 101
rect 1695 648 1745 773
rect 1695 614 1703 648
rect 1737 614 1745 648
rect 1695 580 1745 614
rect 1695 546 1703 580
rect 1737 546 1745 580
rect 1695 512 1745 546
rect 1695 478 1703 512
rect 1737 478 1745 512
rect 1695 185 1745 478
rect 1695 151 1703 185
rect 1737 151 1745 185
rect 1695 67 1745 151
rect 1781 648 1831 773
rect 1781 614 1789 648
rect 1823 614 1831 648
rect 1781 580 1831 614
rect 1781 546 1789 580
rect 1823 546 1831 580
rect 1781 512 1831 546
rect 1781 478 1789 512
rect 1823 478 1831 512
rect 1781 101 1831 478
rect 1781 67 1789 101
rect 1823 67 1831 101
rect 1867 648 1917 773
rect 1867 614 1875 648
rect 1909 614 1917 648
rect 1867 580 1917 614
rect 1867 546 1875 580
rect 1909 546 1917 580
rect 1867 512 1917 546
rect 1867 478 1875 512
rect 1909 478 1917 512
rect 1867 185 1917 478
rect 1867 151 1875 185
rect 1909 151 1917 185
rect 1867 67 1917 151
rect 1953 648 2003 773
rect 1953 614 1961 648
rect 1995 614 2003 648
rect 1953 580 2003 614
rect 1953 546 1961 580
rect 1995 546 2003 580
rect 1953 512 2003 546
rect 1953 478 1961 512
rect 1995 478 2003 512
rect 1953 101 2003 478
rect 1953 67 1961 101
rect 1995 67 2003 101
rect 2039 648 2089 773
rect 2039 614 2047 648
rect 2081 614 2089 648
rect 2039 580 2089 614
rect 2039 546 2047 580
rect 2081 546 2089 580
rect 2039 512 2089 546
rect 2039 478 2047 512
rect 2081 478 2089 512
rect 2039 185 2089 478
rect 2039 151 2047 185
rect 2081 151 2089 185
rect 2039 67 2089 151
rect 2125 648 2175 773
rect 2125 614 2133 648
rect 2167 614 2175 648
rect 2125 580 2175 614
rect 2125 546 2133 580
rect 2167 546 2175 580
rect 2125 512 2175 546
rect 2125 478 2133 512
rect 2167 478 2175 512
rect 2125 101 2175 478
rect 2125 67 2133 101
rect 2167 67 2175 101
rect 2211 648 2261 773
rect 2211 614 2219 648
rect 2253 614 2261 648
rect 2211 580 2261 614
rect 2211 546 2219 580
rect 2253 546 2261 580
rect 2211 512 2261 546
rect 2211 478 2219 512
rect 2253 478 2261 512
rect 2211 185 2261 478
rect 2211 151 2219 185
rect 2253 151 2261 185
rect 2211 67 2261 151
<< viali >>
rect 241 2503 275 2537
rect 413 2503 447 2537
rect 585 2503 619 2537
rect 757 2503 791 2537
rect 929 2503 963 2537
rect 1445 2503 1479 2537
rect 1617 2503 1651 2537
rect 1789 2503 1823 2537
rect 1961 2503 1995 2537
rect 2133 2503 2167 2537
rect 241 2083 275 2117
rect 413 2083 447 2117
rect 585 2083 619 2117
rect 757 2083 791 2117
rect 929 2083 963 2117
rect 1445 2083 1479 2117
rect 1617 2083 1651 2117
rect 1789 2083 1823 2117
rect 1961 2083 1995 2117
rect 2133 2083 2167 2117
rect 155 1327 189 1361
rect 241 1243 275 1277
rect 327 1327 361 1361
rect 413 1243 447 1277
rect 499 1327 533 1361
rect 585 1243 619 1277
rect 671 1327 705 1361
rect 757 1243 791 1277
rect 843 1327 877 1361
rect 929 1243 963 1277
rect 1015 1327 1049 1361
rect 1359 1327 1393 1361
rect 1445 1243 1479 1277
rect 1531 1327 1565 1361
rect 1617 1243 1651 1277
rect 1703 1327 1737 1361
rect 1789 1243 1823 1277
rect 1875 1327 1909 1361
rect 1961 1243 1995 1277
rect 2047 1327 2081 1361
rect 2133 1243 2167 1277
rect 2219 1327 2253 1361
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
rect 1445 907 1479 941
rect 1617 907 1651 941
rect 1789 907 1823 941
rect 1961 907 1995 941
rect 2133 907 2167 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
rect 413 67 447 101
rect 499 151 533 185
rect 585 67 619 101
rect 671 151 705 185
rect 757 67 791 101
rect 843 151 877 185
rect 929 67 963 101
rect 1015 151 1049 185
rect 1359 151 1393 185
rect 1445 67 1479 101
rect 1531 151 1565 185
rect 1617 67 1651 101
rect 1703 151 1737 185
rect 1789 67 1823 101
rect 1875 151 1909 185
rect 1961 67 1995 101
rect 2047 151 2081 185
rect 2133 67 2167 101
rect 2219 151 2253 185
<< metal1 >>
rect 224 2546 980 2548
rect 224 2537 490 2546
rect 224 2503 241 2537
rect 275 2503 413 2537
rect 447 2503 490 2537
rect 224 2494 490 2503
rect 542 2537 980 2546
rect 542 2503 585 2537
rect 619 2503 757 2537
rect 791 2503 929 2537
rect 963 2503 980 2537
rect 542 2494 980 2503
rect 224 2492 980 2494
rect 1428 2546 2184 2548
rect 1428 2537 1866 2546
rect 1428 2503 1445 2537
rect 1479 2503 1617 2537
rect 1651 2503 1789 2537
rect 1823 2503 1866 2537
rect 1428 2494 1866 2503
rect 1918 2537 2184 2546
rect 1918 2503 1961 2537
rect 1995 2503 2133 2537
rect 2167 2503 2184 2537
rect 1918 2494 2184 2503
rect 1428 2492 2184 2494
rect 224 2126 980 2128
rect 224 2117 576 2126
rect 628 2117 980 2126
rect 224 2083 241 2117
rect 275 2083 413 2117
rect 447 2083 576 2117
rect 628 2083 757 2117
rect 791 2083 929 2117
rect 963 2083 980 2117
rect 224 2074 576 2083
rect 628 2074 980 2083
rect 224 2072 980 2074
rect 1428 2126 2184 2128
rect 1428 2117 1780 2126
rect 1832 2117 2184 2126
rect 1428 2083 1445 2117
rect 1479 2083 1617 2117
rect 1651 2083 1780 2117
rect 1832 2083 1961 2117
rect 1995 2083 2133 2117
rect 2167 2083 2184 2117
rect 1428 2074 1780 2083
rect 1832 2074 2184 2083
rect 1428 2072 2184 2074
rect 138 1370 1066 1372
rect 138 1361 490 1370
rect 542 1361 1066 1370
rect 138 1327 155 1361
rect 189 1327 327 1361
rect 361 1327 490 1361
rect 542 1327 671 1361
rect 705 1327 843 1361
rect 877 1327 1015 1361
rect 1049 1327 1066 1361
rect 138 1318 490 1327
rect 542 1318 1066 1327
rect 138 1316 1066 1318
rect 1342 1370 2270 1372
rect 1342 1361 1866 1370
rect 1918 1361 2270 1370
rect 1342 1327 1359 1361
rect 1393 1327 1531 1361
rect 1565 1327 1703 1361
rect 1737 1327 1866 1361
rect 1918 1327 2047 1361
rect 2081 1327 2219 1361
rect 2253 1327 2270 1361
rect 1342 1318 1866 1327
rect 1918 1318 2270 1327
rect 1342 1316 2270 1318
rect 224 1286 980 1288
rect 224 1277 662 1286
rect 224 1243 241 1277
rect 275 1243 413 1277
rect 447 1243 585 1277
rect 619 1243 662 1277
rect 224 1234 662 1243
rect 714 1277 980 1286
rect 714 1243 757 1277
rect 791 1243 929 1277
rect 963 1243 980 1277
rect 714 1234 980 1243
rect 224 1232 980 1234
rect 1428 1286 2184 1288
rect 1428 1277 1694 1286
rect 1428 1243 1445 1277
rect 1479 1243 1617 1277
rect 1651 1243 1694 1277
rect 1428 1234 1694 1243
rect 1746 1277 2184 1286
rect 1746 1243 1789 1277
rect 1823 1243 1961 1277
rect 1995 1243 2133 1277
rect 2167 1243 2184 1277
rect 1746 1234 2184 1243
rect 1428 1232 2184 1234
rect 570 1034 1838 1036
rect 570 982 576 1034
rect 628 982 1780 1034
rect 1832 982 1838 1034
rect 570 980 1838 982
rect 224 950 980 952
rect 224 941 576 950
rect 628 941 980 950
rect 224 907 241 941
rect 275 907 413 941
rect 447 907 576 941
rect 628 907 757 941
rect 791 907 929 941
rect 963 907 980 941
rect 224 898 576 907
rect 628 898 980 907
rect 224 896 980 898
rect 1428 950 2184 952
rect 1428 941 1780 950
rect 1832 941 2184 950
rect 1428 907 1445 941
rect 1479 907 1617 941
rect 1651 907 1780 941
rect 1832 907 1961 941
rect 1995 907 2133 941
rect 2167 907 2184 941
rect 1428 898 1780 907
rect 1832 898 2184 907
rect 1428 896 2184 898
rect 656 278 1752 280
rect 656 226 662 278
rect 714 226 1694 278
rect 1746 226 1752 278
rect 656 224 1752 226
rect 138 194 1066 196
rect 138 185 490 194
rect 542 185 1066 194
rect 138 151 155 185
rect 189 151 327 185
rect 361 151 490 185
rect 542 151 671 185
rect 705 151 843 185
rect 877 151 1015 185
rect 1049 151 1066 185
rect 138 142 490 151
rect 542 142 1066 151
rect 138 140 1066 142
rect 1342 194 2270 196
rect 1342 185 1866 194
rect 1918 185 2270 194
rect 1342 151 1359 185
rect 1393 151 1531 185
rect 1565 151 1703 185
rect 1737 151 1866 185
rect 1918 151 2047 185
rect 2081 151 2219 185
rect 2253 151 2270 185
rect 1342 142 1866 151
rect 1918 142 2270 151
rect 1342 140 2270 142
rect 224 110 980 112
rect 224 101 662 110
rect 224 67 241 101
rect 275 67 413 101
rect 447 67 585 101
rect 619 67 662 101
rect 224 58 662 67
rect 714 101 980 110
rect 714 67 757 101
rect 791 67 929 101
rect 963 67 980 101
rect 714 58 980 67
rect 224 56 980 58
rect 1428 110 2184 112
rect 1428 101 1694 110
rect 1428 67 1445 101
rect 1479 67 1617 101
rect 1651 67 1694 101
rect 1428 58 1694 67
rect 1746 101 2184 110
rect 1746 67 1789 101
rect 1823 67 1961 101
rect 1995 67 2133 101
rect 2167 67 2184 101
rect 1746 58 2184 67
rect 1428 56 2184 58
<< via1 >>
rect 490 2494 542 2546
rect 1866 2494 1918 2546
rect 576 2117 628 2126
rect 576 2083 585 2117
rect 585 2083 619 2117
rect 619 2083 628 2117
rect 576 2074 628 2083
rect 1780 2117 1832 2126
rect 1780 2083 1789 2117
rect 1789 2083 1823 2117
rect 1823 2083 1832 2117
rect 1780 2074 1832 2083
rect 490 1361 542 1370
rect 490 1327 499 1361
rect 499 1327 533 1361
rect 533 1327 542 1361
rect 490 1318 542 1327
rect 1866 1361 1918 1370
rect 1866 1327 1875 1361
rect 1875 1327 1909 1361
rect 1909 1327 1918 1361
rect 1866 1318 1918 1327
rect 662 1234 714 1286
rect 1694 1234 1746 1286
rect 576 982 628 1034
rect 1780 982 1832 1034
rect 576 941 628 950
rect 576 907 585 941
rect 585 907 619 941
rect 619 907 628 941
rect 576 898 628 907
rect 1780 941 1832 950
rect 1780 907 1789 941
rect 1789 907 1823 941
rect 1823 907 1832 941
rect 1780 898 1832 907
rect 662 226 714 278
rect 1694 226 1746 278
rect 490 185 542 194
rect 490 151 499 185
rect 499 151 533 185
rect 533 151 542 185
rect 490 142 542 151
rect 1866 185 1918 194
rect 1866 151 1875 185
rect 1875 151 1909 185
rect 1909 151 1918 185
rect 1866 142 1918 151
rect 662 58 714 110
rect 1694 58 1746 110
<< metal2 >>
rect 488 2546 544 2552
rect 488 2494 490 2546
rect 542 2494 544 2546
rect 488 1370 544 2494
rect 1864 2546 1920 2552
rect 1864 2494 1866 2546
rect 1918 2494 1920 2546
rect 488 1318 490 1370
rect 542 1318 544 1370
rect 488 280 544 1318
rect 574 2126 630 2132
rect 574 2074 576 2126
rect 628 2074 630 2126
rect 574 1034 630 2074
rect 1778 2126 1834 2132
rect 1778 2074 1780 2126
rect 1832 2074 1834 2126
rect 574 982 576 1034
rect 628 982 630 1034
rect 574 950 630 982
rect 574 898 576 950
rect 628 898 630 950
rect 574 892 630 898
rect 660 1286 716 1292
rect 660 1234 662 1286
rect 714 1234 716 1286
rect 488 194 544 224
rect 488 142 490 194
rect 542 142 544 194
rect 488 136 544 142
rect 660 278 716 1234
rect 660 226 662 278
rect 714 226 716 278
rect 660 110 716 226
rect 660 58 662 110
rect 714 58 716 110
rect 660 52 716 58
rect 1692 1286 1748 1292
rect 1692 1234 1694 1286
rect 1746 1234 1748 1286
rect 1692 278 1748 1234
rect 1778 1034 1834 2074
rect 1778 982 1780 1034
rect 1832 982 1834 1034
rect 1778 950 1834 982
rect 1778 898 1780 950
rect 1832 898 1834 950
rect 1778 892 1834 898
rect 1864 1792 1920 2494
rect 1864 1370 1920 1736
rect 1864 1318 1866 1370
rect 1918 1318 1920 1370
rect 1692 226 1694 278
rect 1746 226 1748 278
rect 1692 110 1748 226
rect 1864 194 1920 1318
rect 1864 142 1866 194
rect 1918 142 1920 194
rect 1864 136 1920 142
rect 1692 58 1694 110
rect 1746 58 1748 110
rect 1692 52 1748 58
<< via2 >>
rect 488 224 544 280
rect 1864 1736 1920 1792
<< metal3 >>
rect -80 1796 2448 1844
rect -80 1792 2336 1796
rect -80 1736 1864 1792
rect 1920 1736 2336 1792
rect -80 1732 2336 1736
rect 2400 1732 2448 1796
rect -80 1684 2448 1732
rect 483 284 625 332
rect 483 280 560 284
rect 483 224 488 280
rect 544 224 560 280
rect 483 220 560 224
rect 624 220 625 284
rect 483 172 625 220
rect -80 32 2448 80
rect -80 -32 -32 32
rect 32 -32 560 32
rect 624 -32 2448 32
rect -80 -80 2448 -32
<< via3 >>
rect 2336 1732 2400 1796
rect 560 220 624 284
rect -32 -32 32 32
rect 560 -32 624 32
<< metal4 >>
rect -118 32 118 1882
rect 2250 1796 2486 1882
rect 2250 1732 2336 1796
rect 2400 1732 2486 1796
rect -118 -32 -32 32
rect 32 -32 118 32
rect -118 -118 118 -32
rect 474 284 710 285
rect 474 220 560 284
rect 624 220 710 284
rect 474 32 710 220
rect 474 -32 560 32
rect 624 -32 710 32
rect 474 -33 710 -32
rect 2250 -118 2486 1732
<< labels >>
flabel metal2 s 688 672 688 672 0 FreeSerif 0 0 0 0 Y
port 3 nsew
flabel metal2 s 602 1512 602 1512 0 FreeSerif 0 0 0 0 A
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
port 0 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
port 0 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 1 nsew
flabel metal3 s 554 252 554 252 0 FreeSerif 0 0 0 0 VDD
port 1 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 1 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 1 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 1 nsew
<< end >>
