magic
tech sky130A
magscale 1 2
timestamp 1374899056
<< checkpaint >>
rect -1260 -1260 2464 3948
<< nwell >>
rect 0 0 1204 2688
<< pmos >>
rect 200 1659 230 1827
rect 286 1659 316 1827
rect 372 1659 402 1827
rect 458 1659 488 1827
rect 544 1659 574 1827
rect 630 1659 660 1827
rect 716 1659 746 1827
rect 802 1659 832 1827
rect 888 1659 918 1827
rect 974 1659 1004 1827
rect 200 483 230 651
rect 286 483 316 651
rect 372 483 402 651
rect 458 483 488 651
rect 544 483 574 651
rect 630 483 660 651
rect 716 483 746 651
rect 802 483 832 651
rect 888 483 918 651
rect 974 483 1004 651
<< pdiff >>
rect 147 1777 200 1827
rect 147 1743 155 1777
rect 189 1743 200 1777
rect 147 1709 200 1743
rect 147 1675 155 1709
rect 189 1675 200 1709
rect 147 1659 200 1675
rect 230 1777 286 1827
rect 230 1743 241 1777
rect 275 1743 286 1777
rect 230 1709 286 1743
rect 230 1675 241 1709
rect 275 1675 286 1709
rect 230 1659 286 1675
rect 316 1777 372 1827
rect 316 1743 327 1777
rect 361 1743 372 1777
rect 316 1709 372 1743
rect 316 1675 327 1709
rect 361 1675 372 1709
rect 316 1659 372 1675
rect 402 1777 458 1827
rect 402 1743 413 1777
rect 447 1743 458 1777
rect 402 1709 458 1743
rect 402 1675 413 1709
rect 447 1675 458 1709
rect 402 1659 458 1675
rect 488 1777 544 1827
rect 488 1743 499 1777
rect 533 1743 544 1777
rect 488 1709 544 1743
rect 488 1675 499 1709
rect 533 1675 544 1709
rect 488 1659 544 1675
rect 574 1777 630 1827
rect 574 1743 585 1777
rect 619 1743 630 1777
rect 574 1709 630 1743
rect 574 1675 585 1709
rect 619 1675 630 1709
rect 574 1659 630 1675
rect 660 1777 716 1827
rect 660 1743 671 1777
rect 705 1743 716 1777
rect 660 1709 716 1743
rect 660 1675 671 1709
rect 705 1675 716 1709
rect 660 1659 716 1675
rect 746 1777 802 1827
rect 746 1743 757 1777
rect 791 1743 802 1777
rect 746 1709 802 1743
rect 746 1675 757 1709
rect 791 1675 802 1709
rect 746 1659 802 1675
rect 832 1777 888 1827
rect 832 1743 843 1777
rect 877 1743 888 1777
rect 832 1709 888 1743
rect 832 1675 843 1709
rect 877 1675 888 1709
rect 832 1659 888 1675
rect 918 1777 974 1827
rect 918 1743 929 1777
rect 963 1743 974 1777
rect 918 1709 974 1743
rect 918 1675 929 1709
rect 963 1675 974 1709
rect 918 1659 974 1675
rect 1004 1777 1057 1827
rect 1004 1743 1015 1777
rect 1049 1743 1057 1777
rect 1004 1709 1057 1743
rect 1004 1675 1015 1709
rect 1049 1675 1057 1709
rect 1004 1659 1057 1675
rect 147 601 200 651
rect 147 567 155 601
rect 189 567 200 601
rect 147 533 200 567
rect 147 499 155 533
rect 189 499 200 533
rect 147 483 200 499
rect 230 601 286 651
rect 230 567 241 601
rect 275 567 286 601
rect 230 533 286 567
rect 230 499 241 533
rect 275 499 286 533
rect 230 483 286 499
rect 316 601 372 651
rect 316 567 327 601
rect 361 567 372 601
rect 316 533 372 567
rect 316 499 327 533
rect 361 499 372 533
rect 316 483 372 499
rect 402 601 458 651
rect 402 567 413 601
rect 447 567 458 601
rect 402 533 458 567
rect 402 499 413 533
rect 447 499 458 533
rect 402 483 458 499
rect 488 601 544 651
rect 488 567 499 601
rect 533 567 544 601
rect 488 533 544 567
rect 488 499 499 533
rect 533 499 544 533
rect 488 483 544 499
rect 574 601 630 651
rect 574 567 585 601
rect 619 567 630 601
rect 574 533 630 567
rect 574 499 585 533
rect 619 499 630 533
rect 574 483 630 499
rect 660 601 716 651
rect 660 567 671 601
rect 705 567 716 601
rect 660 533 716 567
rect 660 499 671 533
rect 705 499 716 533
rect 660 483 716 499
rect 746 601 802 651
rect 746 567 757 601
rect 791 567 802 601
rect 746 533 802 567
rect 746 499 757 533
rect 791 499 802 533
rect 746 483 802 499
rect 832 601 888 651
rect 832 567 843 601
rect 877 567 888 601
rect 832 533 888 567
rect 832 499 843 533
rect 877 499 888 533
rect 832 483 888 499
rect 918 601 974 651
rect 918 567 929 601
rect 963 567 974 601
rect 918 533 974 567
rect 918 499 929 533
rect 963 499 974 533
rect 918 483 974 499
rect 1004 601 1057 651
rect 1004 567 1015 601
rect 1049 567 1057 601
rect 1004 533 1057 567
rect 1004 499 1015 533
rect 1049 499 1057 533
rect 1004 483 1057 499
<< pdiffc >>
rect 155 1743 189 1777
rect 155 1675 189 1709
rect 241 1743 275 1777
rect 241 1675 275 1709
rect 327 1743 361 1777
rect 327 1675 361 1709
rect 413 1743 447 1777
rect 413 1675 447 1709
rect 499 1743 533 1777
rect 499 1675 533 1709
rect 585 1743 619 1777
rect 585 1675 619 1709
rect 671 1743 705 1777
rect 671 1675 705 1709
rect 757 1743 791 1777
rect 757 1675 791 1709
rect 843 1743 877 1777
rect 843 1675 877 1709
rect 929 1743 963 1777
rect 929 1675 963 1709
rect 1015 1743 1049 1777
rect 1015 1675 1049 1709
rect 155 567 189 601
rect 155 499 189 533
rect 241 567 275 601
rect 241 499 275 533
rect 327 567 361 601
rect 327 499 361 533
rect 413 567 447 601
rect 413 499 447 533
rect 499 567 533 601
rect 499 499 533 533
rect 585 567 619 601
rect 585 499 619 533
rect 671 567 705 601
rect 671 499 705 533
rect 757 567 791 601
rect 757 499 791 533
rect 843 567 877 601
rect 843 499 877 533
rect 929 567 963 601
rect 929 499 963 533
rect 1015 567 1049 601
rect 1015 499 1049 533
<< nsubdiff >>
rect 241 2537 275 2632
rect 241 2408 275 2503
rect 413 2537 447 2632
rect 413 2408 447 2503
rect 585 2537 619 2632
rect 585 2408 619 2503
rect 757 2537 791 2632
rect 757 2408 791 2503
rect 929 2537 963 2632
rect 929 2408 963 2503
<< nsubdiffcont >>
rect 241 2503 275 2537
rect 413 2503 447 2537
rect 585 2503 619 2537
rect 757 2503 791 2537
rect 929 2503 963 2537
<< poly >>
rect 200 2117 316 2127
rect 200 2083 241 2117
rect 275 2083 316 2117
rect 200 2073 316 2083
rect 200 1827 230 2073
rect 286 1827 316 2073
rect 372 2117 488 2127
rect 372 2083 413 2117
rect 447 2083 488 2117
rect 372 2073 488 2083
rect 372 1827 402 2073
rect 458 1827 488 2073
rect 544 2117 660 2127
rect 544 2083 585 2117
rect 619 2083 660 2117
rect 544 2073 660 2083
rect 544 1827 574 2073
rect 630 1827 660 2073
rect 716 2117 832 2127
rect 716 2083 757 2117
rect 791 2083 832 2117
rect 716 2073 832 2083
rect 716 1827 746 2073
rect 802 1827 832 2073
rect 888 2117 1004 2127
rect 888 2083 929 2117
rect 963 2083 1004 2117
rect 888 2073 1004 2083
rect 888 1827 918 2073
rect 974 1827 1004 2073
rect 200 1428 230 1659
rect 286 1428 316 1659
rect 372 1428 402 1659
rect 458 1428 488 1659
rect 544 1428 574 1659
rect 630 1428 660 1659
rect 716 1428 746 1659
rect 802 1428 832 1659
rect 888 1428 918 1659
rect 974 1428 1004 1659
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 651 230 897
rect 286 651 316 897
rect 372 941 488 951
rect 372 907 413 941
rect 447 907 488 941
rect 372 897 488 907
rect 372 651 402 897
rect 458 651 488 897
rect 544 941 660 951
rect 544 907 585 941
rect 619 907 660 941
rect 544 897 660 907
rect 544 651 574 897
rect 630 651 660 897
rect 716 941 832 951
rect 716 907 757 941
rect 791 907 832 941
rect 716 897 832 907
rect 716 651 746 897
rect 802 651 832 897
rect 888 941 1004 951
rect 888 907 929 941
rect 963 907 1004 941
rect 888 897 1004 907
rect 888 651 918 897
rect 974 651 1004 897
rect 200 252 230 483
rect 286 252 316 483
rect 372 252 402 483
rect 458 252 488 483
rect 544 252 574 483
rect 630 252 660 483
rect 716 252 746 483
rect 802 252 832 483
rect 888 252 918 483
rect 974 252 1004 483
<< polycont >>
rect 241 2083 275 2117
rect 413 2083 447 2117
rect 585 2083 619 2117
rect 757 2083 791 2117
rect 929 2083 963 2117
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
<< locali >>
rect 233 2537 283 2621
rect 233 2503 241 2537
rect 275 2503 283 2537
rect 233 2419 283 2503
rect 405 2537 455 2621
rect 405 2503 413 2537
rect 447 2503 455 2537
rect 405 2419 455 2503
rect 577 2537 627 2621
rect 577 2503 585 2537
rect 619 2503 627 2537
rect 577 2419 627 2503
rect 749 2537 799 2621
rect 749 2503 757 2537
rect 791 2503 799 2537
rect 749 2419 799 2503
rect 921 2537 971 2621
rect 921 2503 929 2537
rect 963 2503 971 2537
rect 921 2419 971 2503
rect 233 2117 283 2201
rect 233 2083 241 2117
rect 275 2083 283 2117
rect 233 1999 283 2083
rect 405 2117 455 2201
rect 405 2083 413 2117
rect 447 2083 455 2117
rect 405 1999 455 2083
rect 577 2117 627 2201
rect 577 2083 585 2117
rect 619 2083 627 2117
rect 577 1999 627 2083
rect 749 2117 799 2201
rect 749 2083 757 2117
rect 791 2083 799 2117
rect 749 1999 799 2083
rect 921 2117 971 2201
rect 921 2083 929 2117
rect 963 2083 971 2117
rect 921 1999 971 2083
rect 147 1777 197 1949
rect 147 1743 155 1777
rect 189 1743 197 1777
rect 147 1709 197 1743
rect 147 1675 155 1709
rect 189 1675 197 1709
rect 147 1361 197 1675
rect 147 1327 155 1361
rect 189 1327 197 1361
rect 147 1243 197 1327
rect 233 1777 283 1949
rect 233 1743 241 1777
rect 275 1743 283 1777
rect 233 1709 283 1743
rect 233 1675 241 1709
rect 275 1675 283 1709
rect 233 1277 283 1675
rect 233 1243 241 1277
rect 275 1243 283 1277
rect 319 1777 369 1949
rect 319 1743 327 1777
rect 361 1743 369 1777
rect 319 1709 369 1743
rect 319 1675 327 1709
rect 361 1675 369 1709
rect 319 1361 369 1675
rect 319 1327 327 1361
rect 361 1327 369 1361
rect 319 1243 369 1327
rect 405 1777 455 1949
rect 405 1743 413 1777
rect 447 1743 455 1777
rect 405 1709 455 1743
rect 405 1675 413 1709
rect 447 1675 455 1709
rect 405 1277 455 1675
rect 405 1243 413 1277
rect 447 1243 455 1277
rect 491 1777 541 1949
rect 491 1743 499 1777
rect 533 1743 541 1777
rect 491 1709 541 1743
rect 491 1675 499 1709
rect 533 1675 541 1709
rect 491 1361 541 1675
rect 491 1327 499 1361
rect 533 1327 541 1361
rect 491 1243 541 1327
rect 577 1777 627 1949
rect 577 1743 585 1777
rect 619 1743 627 1777
rect 577 1709 627 1743
rect 577 1675 585 1709
rect 619 1675 627 1709
rect 577 1277 627 1675
rect 577 1243 585 1277
rect 619 1243 627 1277
rect 663 1777 713 1949
rect 663 1743 671 1777
rect 705 1743 713 1777
rect 663 1709 713 1743
rect 663 1675 671 1709
rect 705 1675 713 1709
rect 663 1361 713 1675
rect 663 1327 671 1361
rect 705 1327 713 1361
rect 663 1243 713 1327
rect 749 1777 799 1949
rect 749 1743 757 1777
rect 791 1743 799 1777
rect 749 1709 799 1743
rect 749 1675 757 1709
rect 791 1675 799 1709
rect 749 1277 799 1675
rect 749 1243 757 1277
rect 791 1243 799 1277
rect 835 1777 885 1949
rect 835 1743 843 1777
rect 877 1743 885 1777
rect 835 1709 885 1743
rect 835 1675 843 1709
rect 877 1675 885 1709
rect 835 1361 885 1675
rect 835 1327 843 1361
rect 877 1327 885 1361
rect 835 1243 885 1327
rect 921 1777 971 1949
rect 921 1743 929 1777
rect 963 1743 971 1777
rect 921 1709 971 1743
rect 921 1675 929 1709
rect 963 1675 971 1709
rect 921 1277 971 1675
rect 921 1243 929 1277
rect 963 1243 971 1277
rect 1007 1777 1057 1949
rect 1007 1743 1015 1777
rect 1049 1743 1057 1777
rect 1007 1709 1057 1743
rect 1007 1675 1015 1709
rect 1049 1675 1057 1709
rect 1007 1361 1057 1675
rect 1007 1327 1015 1361
rect 1049 1327 1057 1361
rect 1007 1243 1057 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 405 941 455 1025
rect 405 907 413 941
rect 447 907 455 941
rect 405 823 455 907
rect 577 941 627 1025
rect 577 907 585 941
rect 619 907 627 941
rect 577 823 627 907
rect 749 941 799 1025
rect 749 907 757 941
rect 791 907 799 941
rect 749 823 799 907
rect 921 941 971 1025
rect 921 907 929 941
rect 963 907 971 941
rect 921 823 971 907
rect 147 601 197 773
rect 147 567 155 601
rect 189 567 197 601
rect 147 533 197 567
rect 147 499 155 533
rect 189 499 197 533
rect 147 185 197 499
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 601 283 773
rect 233 567 241 601
rect 275 567 283 601
rect 233 533 283 567
rect 233 499 241 533
rect 275 499 283 533
rect 233 101 283 499
rect 233 67 241 101
rect 275 67 283 101
rect 319 601 369 773
rect 319 567 327 601
rect 361 567 369 601
rect 319 533 369 567
rect 319 499 327 533
rect 361 499 369 533
rect 319 185 369 499
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
rect 405 601 455 773
rect 405 567 413 601
rect 447 567 455 601
rect 405 533 455 567
rect 405 499 413 533
rect 447 499 455 533
rect 405 101 455 499
rect 405 67 413 101
rect 447 67 455 101
rect 491 601 541 773
rect 491 567 499 601
rect 533 567 541 601
rect 491 533 541 567
rect 491 499 499 533
rect 533 499 541 533
rect 491 185 541 499
rect 491 151 499 185
rect 533 151 541 185
rect 491 67 541 151
rect 577 601 627 773
rect 577 567 585 601
rect 619 567 627 601
rect 577 533 627 567
rect 577 499 585 533
rect 619 499 627 533
rect 577 101 627 499
rect 577 67 585 101
rect 619 67 627 101
rect 663 601 713 773
rect 663 567 671 601
rect 705 567 713 601
rect 663 533 713 567
rect 663 499 671 533
rect 705 499 713 533
rect 663 185 713 499
rect 663 151 671 185
rect 705 151 713 185
rect 663 67 713 151
rect 749 601 799 773
rect 749 567 757 601
rect 791 567 799 601
rect 749 533 799 567
rect 749 499 757 533
rect 791 499 799 533
rect 749 101 799 499
rect 749 67 757 101
rect 791 67 799 101
rect 835 601 885 773
rect 835 567 843 601
rect 877 567 885 601
rect 835 533 885 567
rect 835 499 843 533
rect 877 499 885 533
rect 835 185 885 499
rect 835 151 843 185
rect 877 151 885 185
rect 835 67 885 151
rect 921 601 971 773
rect 921 567 929 601
rect 963 567 971 601
rect 921 533 971 567
rect 921 499 929 533
rect 963 499 971 533
rect 921 101 971 499
rect 921 67 929 101
rect 963 67 971 101
rect 1007 601 1057 773
rect 1007 567 1015 601
rect 1049 567 1057 601
rect 1007 533 1057 567
rect 1007 499 1015 533
rect 1049 499 1057 533
rect 1007 185 1057 499
rect 1007 151 1015 185
rect 1049 151 1057 185
rect 1007 67 1057 151
<< viali >>
rect 241 2503 275 2537
rect 413 2503 447 2537
rect 585 2503 619 2537
rect 757 2503 791 2537
rect 929 2503 963 2537
rect 241 2083 275 2117
rect 413 2083 447 2117
rect 585 2083 619 2117
rect 757 2083 791 2117
rect 929 2083 963 2117
rect 155 1327 189 1361
rect 241 1243 275 1277
rect 327 1327 361 1361
rect 413 1243 447 1277
rect 499 1327 533 1361
rect 585 1243 619 1277
rect 671 1327 705 1361
rect 757 1243 791 1277
rect 843 1327 877 1361
rect 929 1243 963 1277
rect 1015 1327 1049 1361
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
rect 413 67 447 101
rect 499 151 533 185
rect 585 67 619 101
rect 671 151 705 185
rect 757 67 791 101
rect 843 151 877 185
rect 929 67 963 101
rect 1015 151 1049 185
<< metal1 >>
rect 224 2546 980 2548
rect 224 2537 662 2546
rect 224 2503 241 2537
rect 275 2503 413 2537
rect 447 2503 585 2537
rect 619 2503 662 2537
rect 224 2494 662 2503
rect 714 2537 980 2546
rect 714 2503 757 2537
rect 791 2503 929 2537
rect 963 2503 980 2537
rect 714 2494 980 2503
rect 224 2492 980 2494
rect 224 2126 980 2128
rect 224 2117 576 2126
rect 628 2117 980 2126
rect 224 2083 241 2117
rect 275 2083 413 2117
rect 447 2083 576 2117
rect 628 2083 757 2117
rect 791 2083 929 2117
rect 963 2083 980 2117
rect 224 2074 576 2083
rect 628 2074 980 2083
rect 224 2072 980 2074
rect 138 1370 1066 1372
rect 138 1361 662 1370
rect 714 1361 1066 1370
rect 138 1327 155 1361
rect 189 1327 327 1361
rect 361 1327 499 1361
rect 533 1327 662 1361
rect 714 1327 843 1361
rect 877 1327 1015 1361
rect 1049 1327 1066 1361
rect 138 1318 662 1327
rect 714 1318 1066 1327
rect 138 1316 1066 1318
rect 224 1286 980 1288
rect 224 1277 490 1286
rect 224 1243 241 1277
rect 275 1243 413 1277
rect 447 1243 490 1277
rect 224 1234 490 1243
rect 542 1277 980 1286
rect 542 1243 585 1277
rect 619 1243 757 1277
rect 791 1243 929 1277
rect 963 1243 980 1277
rect 542 1234 980 1243
rect 224 1232 980 1234
rect 224 950 980 952
rect 224 941 576 950
rect 628 941 980 950
rect 224 907 241 941
rect 275 907 413 941
rect 447 907 576 941
rect 628 907 757 941
rect 791 907 929 941
rect 963 907 980 941
rect 224 898 576 907
rect 628 898 980 907
rect 224 896 980 898
rect 138 194 1066 196
rect 138 185 662 194
rect 714 185 1066 194
rect 138 151 155 185
rect 189 151 327 185
rect 361 151 499 185
rect 533 151 662 185
rect 714 151 843 185
rect 877 151 1015 185
rect 1049 151 1066 185
rect 138 142 662 151
rect 714 142 1066 151
rect 138 140 1066 142
rect 224 110 980 112
rect 224 101 490 110
rect 224 67 241 101
rect 275 67 413 101
rect 447 67 490 101
rect 224 58 490 67
rect 542 101 980 110
rect 542 67 585 101
rect 619 67 757 101
rect 791 67 929 101
rect 963 67 980 101
rect 542 58 980 67
rect 224 56 980 58
<< via1 >>
rect 662 2494 714 2546
rect 576 2117 628 2126
rect 576 2083 585 2117
rect 585 2083 619 2117
rect 619 2083 628 2117
rect 576 2074 628 2083
rect 662 1361 714 1370
rect 662 1327 671 1361
rect 671 1327 705 1361
rect 705 1327 714 1361
rect 662 1318 714 1327
rect 490 1234 542 1286
rect 576 941 628 950
rect 576 907 585 941
rect 585 907 619 941
rect 619 907 628 941
rect 576 898 628 907
rect 662 185 714 194
rect 662 151 671 185
rect 671 151 705 185
rect 705 151 714 185
rect 662 142 714 151
rect 490 58 542 110
<< metal2 >>
rect 660 2546 716 2552
rect 660 2494 662 2546
rect 714 2494 716 2546
rect 574 2126 630 2132
rect 574 2074 576 2126
rect 628 2074 630 2126
rect 488 1286 544 1292
rect 488 1234 490 1286
rect 542 1234 544 1286
rect 488 110 544 1234
rect 574 950 630 2074
rect 574 898 576 950
rect 628 898 630 950
rect 574 892 630 898
rect 660 1370 716 2494
rect 660 1318 662 1370
rect 714 1318 716 1370
rect 660 194 716 1318
rect 660 142 662 194
rect 714 142 716 194
rect 660 136 716 142
rect 488 58 490 110
rect 542 58 544 110
rect 488 52 544 58
<< end >>
