magic
tech sky130A
magscale 1 2
timestamp 1614649966
<< nwell >>
rect -110 247 2082 568
<< pwell >>
rect -43 50 -9 155
rect 1981 50 2015 155
rect 49 -31 83 3
rect 325 -31 359 3
rect 601 -31 635 3
rect 877 -31 911 3
rect 1153 -31 1187 3
rect 1429 -31 1463 3
rect 1705 -31 1739 3
<< scnmos >>
rect 140 33 170 163
rect 416 33 446 163
rect 692 33 722 163
rect 968 33 998 163
rect 1244 33 1274 163
rect 1520 33 1550 163
rect 1796 33 1826 163
<< scpmoshvt >>
rect 140 283 170 483
rect 416 283 446 483
rect 692 283 722 483
rect 968 283 998 483
rect 1244 283 1274 483
rect 1520 283 1550 483
rect 1796 283 1826 483
<< ndiff >>
rect 88 151 140 163
rect 88 117 96 151
rect 130 117 140 151
rect 88 83 140 117
rect 88 49 96 83
rect 130 49 140 83
rect 88 33 140 49
rect 170 151 222 163
rect 170 117 180 151
rect 214 117 222 151
rect 170 83 222 117
rect 170 49 180 83
rect 214 49 222 83
rect 170 33 222 49
rect 364 151 416 163
rect 364 117 372 151
rect 406 117 416 151
rect 364 83 416 117
rect 364 49 372 83
rect 406 49 416 83
rect 364 33 416 49
rect 446 151 498 163
rect 446 117 456 151
rect 490 117 498 151
rect 446 83 498 117
rect 446 49 456 83
rect 490 49 498 83
rect 446 33 498 49
rect 640 151 692 163
rect 640 117 648 151
rect 682 117 692 151
rect 640 83 692 117
rect 640 49 648 83
rect 682 49 692 83
rect 640 33 692 49
rect 722 151 774 163
rect 722 117 732 151
rect 766 117 774 151
rect 722 83 774 117
rect 722 49 732 83
rect 766 49 774 83
rect 722 33 774 49
rect 916 151 968 163
rect 916 117 924 151
rect 958 117 968 151
rect 916 83 968 117
rect 916 49 924 83
rect 958 49 968 83
rect 916 33 968 49
rect 998 151 1050 163
rect 998 117 1008 151
rect 1042 117 1050 151
rect 998 83 1050 117
rect 998 49 1008 83
rect 1042 49 1050 83
rect 998 33 1050 49
rect 1192 151 1244 163
rect 1192 117 1200 151
rect 1234 117 1244 151
rect 1192 83 1244 117
rect 1192 49 1200 83
rect 1234 49 1244 83
rect 1192 33 1244 49
rect 1274 151 1326 163
rect 1274 117 1284 151
rect 1318 117 1326 151
rect 1274 83 1326 117
rect 1274 49 1284 83
rect 1318 49 1326 83
rect 1274 33 1326 49
rect 1468 151 1520 163
rect 1468 117 1476 151
rect 1510 117 1520 151
rect 1468 83 1520 117
rect 1468 49 1476 83
rect 1510 49 1520 83
rect 1468 33 1520 49
rect 1550 151 1602 163
rect 1550 117 1560 151
rect 1594 117 1602 151
rect 1550 83 1602 117
rect 1550 49 1560 83
rect 1594 49 1602 83
rect 1550 33 1602 49
rect 1744 151 1796 163
rect 1744 117 1752 151
rect 1786 117 1796 151
rect 1744 83 1796 117
rect 1744 49 1752 83
rect 1786 49 1796 83
rect 1744 33 1796 49
rect 1826 151 1878 163
rect 1826 117 1836 151
rect 1870 117 1878 151
rect 1826 83 1878 117
rect 1826 49 1836 83
rect 1870 49 1878 83
rect 1826 33 1878 49
<< pdiff >>
rect 88 471 140 483
rect 88 437 96 471
rect 130 437 140 471
rect 88 403 140 437
rect 88 369 96 403
rect 130 369 140 403
rect 88 335 140 369
rect 88 301 96 335
rect 130 301 140 335
rect 88 283 140 301
rect 170 471 222 483
rect 170 437 180 471
rect 214 437 222 471
rect 170 403 222 437
rect 170 369 180 403
rect 214 369 222 403
rect 170 335 222 369
rect 170 301 180 335
rect 214 301 222 335
rect 170 283 222 301
rect 364 471 416 483
rect 364 437 372 471
rect 406 437 416 471
rect 364 403 416 437
rect 364 369 372 403
rect 406 369 416 403
rect 364 335 416 369
rect 364 301 372 335
rect 406 301 416 335
rect 364 283 416 301
rect 446 471 498 483
rect 446 437 456 471
rect 490 437 498 471
rect 446 403 498 437
rect 446 369 456 403
rect 490 369 498 403
rect 446 335 498 369
rect 446 301 456 335
rect 490 301 498 335
rect 446 283 498 301
rect 640 471 692 483
rect 640 437 648 471
rect 682 437 692 471
rect 640 403 692 437
rect 640 369 648 403
rect 682 369 692 403
rect 640 335 692 369
rect 640 301 648 335
rect 682 301 692 335
rect 640 283 692 301
rect 722 471 774 483
rect 722 437 732 471
rect 766 437 774 471
rect 722 403 774 437
rect 722 369 732 403
rect 766 369 774 403
rect 722 335 774 369
rect 722 301 732 335
rect 766 301 774 335
rect 722 283 774 301
rect 916 471 968 483
rect 916 437 924 471
rect 958 437 968 471
rect 916 403 968 437
rect 916 369 924 403
rect 958 369 968 403
rect 916 335 968 369
rect 916 301 924 335
rect 958 301 968 335
rect 916 283 968 301
rect 998 471 1050 483
rect 998 437 1008 471
rect 1042 437 1050 471
rect 998 403 1050 437
rect 998 369 1008 403
rect 1042 369 1050 403
rect 998 335 1050 369
rect 998 301 1008 335
rect 1042 301 1050 335
rect 998 283 1050 301
rect 1192 471 1244 483
rect 1192 437 1200 471
rect 1234 437 1244 471
rect 1192 403 1244 437
rect 1192 369 1200 403
rect 1234 369 1244 403
rect 1192 335 1244 369
rect 1192 301 1200 335
rect 1234 301 1244 335
rect 1192 283 1244 301
rect 1274 471 1326 483
rect 1274 437 1284 471
rect 1318 437 1326 471
rect 1274 403 1326 437
rect 1274 369 1284 403
rect 1318 369 1326 403
rect 1274 335 1326 369
rect 1274 301 1284 335
rect 1318 301 1326 335
rect 1274 283 1326 301
rect 1468 471 1520 483
rect 1468 437 1476 471
rect 1510 437 1520 471
rect 1468 403 1520 437
rect 1468 369 1476 403
rect 1510 369 1520 403
rect 1468 335 1520 369
rect 1468 301 1476 335
rect 1510 301 1520 335
rect 1468 283 1520 301
rect 1550 471 1602 483
rect 1550 437 1560 471
rect 1594 437 1602 471
rect 1550 403 1602 437
rect 1550 369 1560 403
rect 1594 369 1602 403
rect 1550 335 1602 369
rect 1550 301 1560 335
rect 1594 301 1602 335
rect 1550 283 1602 301
rect 1744 471 1796 483
rect 1744 437 1752 471
rect 1786 437 1796 471
rect 1744 403 1796 437
rect 1744 369 1752 403
rect 1786 369 1796 403
rect 1744 335 1796 369
rect 1744 301 1752 335
rect 1786 301 1796 335
rect 1744 283 1796 301
rect 1826 471 1878 483
rect 1826 437 1836 471
rect 1870 437 1878 471
rect 1826 403 1878 437
rect 1826 369 1836 403
rect 1870 369 1878 403
rect 1826 335 1878 369
rect 1826 301 1836 335
rect 1870 301 1878 335
rect 1826 283 1878 301
<< ndiffc >>
rect 96 117 130 151
rect 96 49 130 83
rect 180 117 214 151
rect 180 49 214 83
rect 372 117 406 151
rect 372 49 406 83
rect 456 117 490 151
rect 456 49 490 83
rect 648 117 682 151
rect 648 49 682 83
rect 732 117 766 151
rect 732 49 766 83
rect 924 117 958 151
rect 924 49 958 83
rect 1008 117 1042 151
rect 1008 49 1042 83
rect 1200 117 1234 151
rect 1200 49 1234 83
rect 1284 117 1318 151
rect 1284 49 1318 83
rect 1476 117 1510 151
rect 1476 49 1510 83
rect 1560 117 1594 151
rect 1560 49 1594 83
rect 1752 117 1786 151
rect 1752 49 1786 83
rect 1836 117 1870 151
rect 1836 49 1870 83
<< pdiffc >>
rect 96 437 130 471
rect 96 369 130 403
rect 96 301 130 335
rect 180 437 214 471
rect 180 369 214 403
rect 180 301 214 335
rect 372 437 406 471
rect 372 369 406 403
rect 372 301 406 335
rect 456 437 490 471
rect 456 369 490 403
rect 456 301 490 335
rect 648 437 682 471
rect 648 369 682 403
rect 648 301 682 335
rect 732 437 766 471
rect 732 369 766 403
rect 732 301 766 335
rect 924 437 958 471
rect 924 369 958 403
rect 924 301 958 335
rect 1008 437 1042 471
rect 1008 369 1042 403
rect 1008 301 1042 335
rect 1200 437 1234 471
rect 1200 369 1234 403
rect 1200 301 1234 335
rect 1284 437 1318 471
rect 1284 369 1318 403
rect 1284 301 1318 335
rect 1476 437 1510 471
rect 1476 369 1510 403
rect 1476 301 1510 335
rect 1560 437 1594 471
rect 1560 369 1594 403
rect 1560 301 1594 335
rect 1752 437 1786 471
rect 1752 369 1786 403
rect 1752 301 1786 335
rect 1836 437 1870 471
rect 1836 369 1870 403
rect 1836 301 1870 335
<< psubdiff >>
rect -43 131 -9 155
rect -43 50 -9 97
rect 1981 131 2015 155
rect 1981 50 2015 97
<< nsubdiff >>
rect -43 442 -9 466
rect -43 349 -9 408
rect -43 291 -9 315
rect 1981 442 2015 466
rect 1981 349 2015 408
rect 1981 291 2015 315
<< psubdiffcont >>
rect -43 97 -9 131
rect 1981 97 2015 131
<< nsubdiffcont >>
rect -43 408 -9 442
rect -43 315 -9 349
rect 1981 408 2015 442
rect 1981 315 2015 349
<< poly >>
rect 140 483 170 509
rect 416 483 446 509
rect 692 483 722 509
rect 968 483 998 509
rect 1244 483 1274 509
rect 1520 483 1550 509
rect 1796 483 1826 509
rect 140 251 170 283
rect 416 251 446 283
rect 692 251 722 283
rect 968 251 998 283
rect 1244 251 1274 283
rect 1520 251 1550 283
rect 1796 251 1826 283
rect 84 235 170 251
rect 84 201 100 235
rect 134 201 170 235
rect 84 185 170 201
rect 360 235 446 251
rect 360 201 376 235
rect 410 201 446 235
rect 360 185 446 201
rect 636 235 722 251
rect 636 201 652 235
rect 686 201 722 235
rect 636 185 722 201
rect 912 235 998 251
rect 912 201 928 235
rect 962 201 998 235
rect 912 185 998 201
rect 1188 235 1274 251
rect 1188 201 1204 235
rect 1238 201 1274 235
rect 1188 185 1274 201
rect 1464 235 1550 251
rect 1464 201 1480 235
rect 1514 201 1550 235
rect 1464 185 1550 201
rect 1740 235 1826 251
rect 1740 201 1756 235
rect 1790 201 1826 235
rect 1740 185 1826 201
rect 140 163 170 185
rect 416 163 446 185
rect 692 163 722 185
rect 968 163 998 185
rect 1244 163 1274 185
rect 1520 163 1550 185
rect 1796 163 1826 185
rect 140 7 170 33
rect 416 7 446 33
rect 692 7 722 33
rect 968 7 998 33
rect 1244 7 1274 33
rect 1520 7 1550 33
rect 1796 7 1826 33
<< polycont >>
rect 100 201 134 235
rect 376 201 410 235
rect 652 201 686 235
rect 928 201 962 235
rect 1204 201 1238 235
rect 1480 201 1514 235
rect 1756 201 1790 235
<< locali >>
rect -72 513 -43 547
rect -9 513 49 547
rect 83 513 141 547
rect 175 513 233 547
rect 267 513 325 547
rect 359 513 417 547
rect 451 513 509 547
rect 543 513 601 547
rect 635 513 693 547
rect 727 513 785 547
rect 819 513 877 547
rect 911 513 969 547
rect 1003 513 1061 547
rect 1095 513 1153 547
rect 1187 513 1245 547
rect 1279 513 1337 547
rect 1371 513 1429 547
rect 1463 513 1521 547
rect 1555 513 1613 547
rect 1647 513 1705 547
rect 1739 513 1797 547
rect 1831 513 1889 547
rect 1923 513 1981 547
rect 2015 513 2044 547
rect -55 442 3 513
rect -55 408 -43 442
rect -9 408 3 442
rect -55 349 3 408
rect -55 315 -43 349
rect -9 315 3 349
rect -55 280 3 315
rect 88 471 130 513
rect 88 437 96 471
rect 88 403 130 437
rect 88 369 96 403
rect 88 335 130 369
rect 88 301 96 335
rect 88 285 130 301
rect 164 471 230 479
rect 164 437 180 471
rect 214 437 230 471
rect 164 403 230 437
rect 164 369 180 403
rect 214 369 230 403
rect 164 335 230 369
rect 164 301 180 335
rect 214 301 230 335
rect 164 283 230 301
rect 364 471 406 513
rect 364 437 372 471
rect 364 403 406 437
rect 364 369 372 403
rect 364 335 406 369
rect 364 301 372 335
rect 364 285 406 301
rect 440 471 506 479
rect 440 437 456 471
rect 490 437 506 471
rect 440 403 506 437
rect 440 369 456 403
rect 490 369 506 403
rect 440 335 506 369
rect 440 301 456 335
rect 490 301 506 335
rect 440 283 506 301
rect 640 471 682 513
rect 640 437 648 471
rect 640 403 682 437
rect 640 369 648 403
rect 640 335 682 369
rect 640 301 648 335
rect 640 285 682 301
rect 716 471 782 479
rect 716 437 732 471
rect 766 437 782 471
rect 716 403 782 437
rect 716 369 732 403
rect 766 369 782 403
rect 716 335 782 369
rect 716 301 732 335
rect 766 301 782 335
rect 716 283 782 301
rect 916 471 958 513
rect 916 437 924 471
rect 916 403 958 437
rect 916 369 924 403
rect 916 335 958 369
rect 916 301 924 335
rect 916 285 958 301
rect 992 471 1058 479
rect 992 437 1008 471
rect 1042 437 1058 471
rect 992 403 1058 437
rect 992 369 1008 403
rect 1042 369 1058 403
rect 992 335 1058 369
rect 992 301 1008 335
rect 1042 301 1058 335
rect 992 283 1058 301
rect 1192 471 1234 513
rect 1192 437 1200 471
rect 1192 403 1234 437
rect 1192 369 1200 403
rect 1192 335 1234 369
rect 1192 301 1200 335
rect 1192 285 1234 301
rect 1268 471 1334 479
rect 1268 437 1284 471
rect 1318 437 1334 471
rect 1268 403 1334 437
rect 1268 369 1284 403
rect 1318 369 1334 403
rect 1268 335 1334 369
rect 1268 301 1284 335
rect 1318 301 1334 335
rect 1268 283 1334 301
rect 1468 471 1510 513
rect 1468 437 1476 471
rect 1468 403 1510 437
rect 1468 369 1476 403
rect 1468 335 1510 369
rect 1468 301 1476 335
rect 1468 285 1510 301
rect 1544 471 1610 479
rect 1544 437 1560 471
rect 1594 437 1610 471
rect 1544 403 1610 437
rect 1544 369 1560 403
rect 1594 369 1610 403
rect 1544 335 1610 369
rect 1544 301 1560 335
rect 1594 301 1610 335
rect 1544 283 1610 301
rect 1744 471 1786 513
rect 1744 437 1752 471
rect 1744 403 1786 437
rect 1744 369 1752 403
rect 1744 335 1786 369
rect 1744 301 1752 335
rect 1744 285 1786 301
rect 1820 471 1886 479
rect 1820 437 1836 471
rect 1870 437 1886 471
rect 1820 403 1886 437
rect 1820 369 1836 403
rect 1870 369 1886 403
rect 1820 335 1886 369
rect 1820 301 1836 335
rect 1870 301 1886 335
rect 1820 283 1886 301
rect 184 249 230 283
rect 460 249 506 283
rect 736 249 782 283
rect 1012 249 1058 283
rect 1288 249 1334 283
rect 1564 249 1610 283
rect 84 241 150 249
rect 84 207 91 241
rect 125 235 150 241
rect 84 201 100 207
rect 134 201 150 235
rect 184 235 426 249
rect 184 201 376 235
rect 410 201 426 235
rect 460 235 702 249
rect 460 201 652 235
rect 686 201 702 235
rect 736 235 978 249
rect 736 201 928 235
rect 962 201 978 235
rect 1012 235 1254 249
rect 1012 201 1204 235
rect 1238 201 1254 235
rect 1288 235 1530 249
rect 1288 201 1480 235
rect 1514 201 1530 235
rect 1564 235 1806 249
rect 1564 202 1756 235
rect 84 151 130 167
rect 184 163 230 201
rect -55 131 3 148
rect -55 97 -43 131
rect -9 97 3 131
rect -55 3 3 97
rect 84 117 96 151
rect 84 83 130 117
rect 84 49 96 83
rect 84 3 130 49
rect 164 151 230 163
rect 164 117 180 151
rect 214 117 230 151
rect 164 83 230 117
rect 164 49 180 83
rect 214 49 230 83
rect 164 37 230 49
rect 360 151 406 167
rect 460 163 506 201
rect 360 117 372 151
rect 360 83 406 117
rect 360 49 372 83
rect 360 3 406 49
rect 440 151 506 163
rect 440 117 456 151
rect 490 117 506 151
rect 440 83 506 117
rect 440 49 456 83
rect 490 49 506 83
rect 440 37 506 49
rect 636 151 682 167
rect 736 163 782 201
rect 636 117 648 151
rect 636 83 682 117
rect 636 49 648 83
rect 636 3 682 49
rect 716 151 782 163
rect 716 117 732 151
rect 766 117 782 151
rect 716 83 782 117
rect 716 49 732 83
rect 766 49 782 83
rect 716 37 782 49
rect 912 151 958 167
rect 1012 163 1058 201
rect 912 117 924 151
rect 912 83 958 117
rect 912 49 924 83
rect 912 3 958 49
rect 992 151 1058 163
rect 992 117 1008 151
rect 1042 117 1058 151
rect 992 83 1058 117
rect 992 49 1008 83
rect 1042 49 1058 83
rect 992 37 1058 49
rect 1188 151 1234 167
rect 1288 163 1334 201
rect 1188 117 1200 151
rect 1188 83 1234 117
rect 1188 49 1200 83
rect 1188 3 1234 49
rect 1268 151 1334 163
rect 1268 117 1284 151
rect 1318 117 1334 151
rect 1268 83 1334 117
rect 1268 49 1284 83
rect 1318 49 1334 83
rect 1268 37 1334 49
rect 1464 151 1510 167
rect 1564 163 1610 202
rect 1740 201 1756 202
rect 1790 201 1806 235
rect 1840 244 1886 283
rect 1969 442 2027 513
rect 1969 408 1981 442
rect 2015 408 2027 442
rect 1969 349 2027 408
rect 1969 315 1981 349
rect 2015 315 2027 349
rect 1969 280 2027 315
rect 1840 241 2083 244
rect 1840 207 1846 241
rect 1880 207 2083 241
rect 1840 196 2083 207
rect 1464 117 1476 151
rect 1464 83 1510 117
rect 1464 49 1476 83
rect 1464 3 1510 49
rect 1544 151 1610 163
rect 1544 117 1560 151
rect 1594 117 1610 151
rect 1544 83 1610 117
rect 1544 49 1560 83
rect 1594 49 1610 83
rect 1544 37 1610 49
rect 1740 151 1786 167
rect 1840 163 1886 196
rect 1740 117 1752 151
rect 1740 83 1786 117
rect 1740 49 1752 83
rect 1740 3 1786 49
rect 1820 151 1886 163
rect 1820 117 1836 151
rect 1870 117 1886 151
rect 1820 83 1886 117
rect 1820 49 1836 83
rect 1870 49 1886 83
rect 1820 37 1886 49
rect 1969 131 2027 148
rect 1969 97 1981 131
rect 2015 97 2027 131
rect 1969 3 2027 97
rect -72 -31 -43 3
rect -9 -31 49 3
rect 83 -31 141 3
rect 175 -31 233 3
rect 267 -31 325 3
rect 359 -31 417 3
rect 451 -31 509 3
rect 543 -31 601 3
rect 635 -31 693 3
rect 727 -31 785 3
rect 819 -31 877 3
rect 911 -31 969 3
rect 1003 -31 1061 3
rect 1095 -31 1153 3
rect 1187 -31 1245 3
rect 1279 -31 1337 3
rect 1371 -31 1429 3
rect 1463 -31 1521 3
rect 1555 -31 1613 3
rect 1647 -31 1705 3
rect 1739 -31 1797 3
rect 1831 -31 1889 3
rect 1923 -31 1981 3
rect 2015 -31 2044 3
<< viali >>
rect -43 513 -9 547
rect 49 513 83 547
rect 141 513 175 547
rect 233 513 267 547
rect 325 513 359 547
rect 417 513 451 547
rect 509 513 543 547
rect 601 513 635 547
rect 693 513 727 547
rect 785 513 819 547
rect 877 513 911 547
rect 969 513 1003 547
rect 1061 513 1095 547
rect 1153 513 1187 547
rect 1245 513 1279 547
rect 1337 513 1371 547
rect 1429 513 1463 547
rect 1521 513 1555 547
rect 1613 513 1647 547
rect 1705 513 1739 547
rect 1797 513 1831 547
rect 1889 513 1923 547
rect 1981 513 2015 547
rect 91 235 125 241
rect 91 207 100 235
rect 100 207 125 235
rect 1846 207 1880 241
rect -43 -31 -9 3
rect 49 -31 83 3
rect 141 -31 175 3
rect 233 -31 267 3
rect 325 -31 359 3
rect 417 -31 451 3
rect 509 -31 543 3
rect 601 -31 635 3
rect 693 -31 727 3
rect 785 -31 819 3
rect 877 -31 911 3
rect 969 -31 1003 3
rect 1061 -31 1095 3
rect 1153 -31 1187 3
rect 1245 -31 1279 3
rect 1337 -31 1371 3
rect 1429 -31 1463 3
rect 1521 -31 1555 3
rect 1613 -31 1647 3
rect 1705 -31 1739 3
rect 1797 -31 1831 3
rect 1889 -31 1923 3
rect 1981 -31 2015 3
<< metal1 >>
rect -72 547 2082 578
rect -72 513 -43 547
rect -9 513 49 547
rect 83 513 141 547
rect 175 513 233 547
rect 267 513 325 547
rect 359 513 417 547
rect 451 513 509 547
rect 543 513 601 547
rect 635 513 693 547
rect 727 513 785 547
rect 819 513 877 547
rect 911 513 969 547
rect 1003 513 1061 547
rect 1095 513 1153 547
rect 1187 513 1245 547
rect 1279 513 1337 547
rect 1371 513 1429 547
rect 1463 513 1521 547
rect 1555 513 1613 547
rect 1647 513 1705 547
rect 1739 513 1797 547
rect 1831 513 1889 547
rect 1923 513 1981 547
rect 2015 513 2082 547
rect -72 482 2082 513
rect 79 241 1892 253
rect 79 207 91 241
rect 125 207 1846 241
rect 1880 207 1892 241
rect 79 195 1892 207
rect -72 3 2082 34
rect -72 -31 -43 3
rect -9 -31 49 3
rect 83 -31 141 3
rect 175 -31 233 3
rect 267 -31 325 3
rect 359 -31 417 3
rect 451 -31 509 3
rect 543 -31 601 3
rect 635 -31 693 3
rect 727 -31 785 3
rect 819 -31 877 3
rect 911 -31 969 3
rect 1003 -31 1061 3
rect 1095 -31 1153 3
rect 1187 -31 1245 3
rect 1279 -31 1337 3
rect 1371 -31 1429 3
rect 1463 -31 1521 3
rect 1555 -31 1613 3
rect 1647 -31 1705 3
rect 1739 -31 1797 3
rect 1831 -31 1889 3
rect 1923 -31 1981 3
rect 2015 -31 2082 3
rect -72 -62 2082 -31
<< labels >>
flabel locali 1841 196 2083 244 1 FreeSans 400 0 0 0 out
port 1 n
flabel metal1 2044 482 2082 578 1 FreeSans 400 0 0 0 vdd
port 2 n
flabel metal1 2044 -62 2082 34 1 FreeSans 400 0 0 0 gnd
port 3 n
flabel metal1 1974 510 2027 539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 1973 -32 2024 6 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment 1952 -14 1952 -14 4 sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
flabel metal1 -50 510 3 539 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 -51 -32 0 6 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment -72 -14 -72 -14 4 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
flabel locali 184 275 218 309 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[0]/Y
flabel locali 184 207 218 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[0]/Y
flabel locali 92 207 126 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[0]/A
flabel nwell 49 513 83 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[0]/VPB
flabel pwell 49 -31 83 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[0]/VNB
flabel metal1 49 -31 83 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[0]/VGND
flabel metal1 49 513 83 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[0]/VPWR
rlabel comment 20 -14 20 -14 4 sky130_fd_sc_hd__inv_1_0[0]/inv_1
flabel locali 460 275 494 309 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[1]/Y
flabel locali 460 207 494 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[1]/Y
flabel locali 368 207 402 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[1]/A
flabel nwell 325 513 359 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[1]/VPB
flabel pwell 325 -31 359 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[1]/VNB
flabel metal1 325 -31 359 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[1]/VGND
flabel metal1 325 513 359 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[1]/VPWR
rlabel comment 296 -14 296 -14 4 sky130_fd_sc_hd__inv_1_0[1]/inv_1
flabel locali 736 275 770 309 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[2]/Y
flabel locali 736 207 770 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[2]/Y
flabel locali 644 207 678 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[2]/A
flabel nwell 601 513 635 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[2]/VPB
flabel pwell 601 -31 635 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[2]/VNB
flabel metal1 601 -31 635 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[2]/VGND
flabel metal1 601 513 635 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[2]/VPWR
rlabel comment 572 -14 572 -14 4 sky130_fd_sc_hd__inv_1_0[2]/inv_1
flabel locali 1012 275 1046 309 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[3]/Y
flabel locali 1012 207 1046 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[3]/Y
flabel locali 920 207 954 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[3]/A
flabel nwell 877 513 911 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[3]/VPB
flabel pwell 877 -31 911 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[3]/VNB
flabel metal1 877 -31 911 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[3]/VGND
flabel metal1 877 513 911 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[3]/VPWR
rlabel comment 848 -14 848 -14 4 sky130_fd_sc_hd__inv_1_0[3]/inv_1
flabel locali 1288 275 1322 309 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[4]/Y
flabel locali 1288 207 1322 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[4]/Y
flabel locali 1196 207 1230 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[4]/A
flabel nwell 1153 513 1187 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[4]/VPB
flabel pwell 1153 -31 1187 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[4]/VNB
flabel metal1 1153 -31 1187 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[4]/VGND
flabel metal1 1153 513 1187 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[4]/VPWR
rlabel comment 1124 -14 1124 -14 4 sky130_fd_sc_hd__inv_1_0[4]/inv_1
flabel locali 1564 275 1598 309 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[5]/Y
flabel locali 1564 207 1598 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[5]/Y
flabel locali 1472 207 1506 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[5]/A
flabel nwell 1429 513 1463 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[5]/VPB
flabel pwell 1429 -31 1463 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[5]/VNB
flabel metal1 1429 -31 1463 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[5]/VGND
flabel metal1 1429 513 1463 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[5]/VPWR
rlabel comment 1400 -14 1400 -14 4 sky130_fd_sc_hd__inv_1_0[5]/inv_1
flabel locali 1840 275 1874 309 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[6]/Y
flabel locali 1840 207 1874 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[6]/Y
flabel locali 1748 207 1782 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0[6]/A
flabel nwell 1705 513 1739 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[6]/VPB
flabel pwell 1705 -31 1739 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[6]/VNB
flabel metal1 1705 -31 1739 3 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[6]/VGND
flabel metal1 1705 513 1739 547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0[6]/VPWR
rlabel comment 1676 -14 1676 -14 4 sky130_fd_sc_hd__inv_1_0[6]/inv_1
<< end >>
