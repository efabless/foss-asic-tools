* NGSPICE file created from schmittbuf.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__schmittbuf_1 A VGND VNB VPB VPWR X
X0 a_64_207# VPWR VPB sky130_fd_pr__res_generic_pd w=290000u l=3.11e+06u
X1 a_231_463# A a_117_181# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=4.0875e+11p pd=4.09e+06u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X2 a_217_207# A a_117_181# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=2.289e+11p pd=2.77e+06u as=1.113e+11p ps=1.37e+06u w=420000u l=500000u
X3 VPWR A a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=1.02225e+12p pd=5.2e+06u as=0p ps=0u w=750000u l=500000u
X4 a_217_207# a_117_181# a_64_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=500000u
X5 X a_117_181# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=9.478e+11p ps=4.36e+06u w=750000u l=500000u
X6 a_78_463# VGND VNB sky130_fd_pr__res_generic_nd w=290000u l=1.355e+06u
X7 X a_117_181# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X8 VGND A a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X9 a_231_463# a_117_181# a_78_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
C0 VGND A 0.04fF
C1 a_117_181# a_64_207# 0.06fF
C2 VPWR A 0.07fF
C3 a_231_463# a_117_181# 0.32fF
C4 a_78_463# a_117_181# 0.40fF
C5 VPWR a_64_207# 0.13fF
C6 VPWR a_231_463# 0.10fF
C7 a_78_463# VGND 0.15fF
C8 a_217_207# a_117_181# 0.31fF
C9 VPB a_117_181# 0.03fF
C10 a_231_463# A 0.18fF
C11 X VPB 0.05fF
C12 VGND a_217_207# 0.03fF
C13 VPWR VPB 1.91fF
C14 a_231_463# a_64_207# 0.04fF
C15 a_78_463# a_64_207# 0.40fF
C16 a_231_463# a_78_463# 0.07fF
C17 A a_217_207# 0.12fF
C18 A VPB 0.02fF
C19 a_217_207# a_64_207# 0.02fF
C20 VPB a_64_207# 0.12fF
C21 a_231_463# a_217_207# 0.02fF
C22 a_231_463# VPB 0.11fF
C23 a_78_463# a_217_207# 0.26fF
C24 a_78_463# VPB 0.01fF
C25 X a_117_181# 0.28fF
C26 VGND a_117_181# 0.35fF
C27 VGND X 0.16fF
C28 VPWR a_117_181# 0.32fF
C29 VPWR X 0.23fF
C30 VPWR VGND 0.04fF
C31 A a_117_181# 0.57fF
C32 VGND VNB 0.44fF
C33 X VNB 0.22fF
C34 A VNB 0.49fF
C35 VPWR VNB 0.40fF
C36 VPB VNB 2.88fF
C37 a_217_207# VNB 0.13fF
C38 a_231_463# VNB 0.24fF
C39 a_78_463# VNB 0.19fF
C40 a_64_207# VNB 0.41fF
C41 a_117_181# VNB 0.94fF
.ends


* Top level circuit schmittbuf

Xsky130_fd_sc_hvl__schmittbuf_1_0 sky130_fd_sc_hvl__schmittbuf_1_0/A sky130_fd_sc_hvl__schmittbuf_1_0/VGND
+ VSUBS sky130_fd_sc_hvl__schmittbuf_1_0/VPB sky130_fd_sc_hvl__schmittbuf_1_0/VPWR
+ sky130_fd_sc_hvl__schmittbuf_1_0/X sky130_fd_sc_hvl__schmittbuf_1
C0 sky130_fd_sc_hvl__schmittbuf_1_0/VGND VSUBS 0.44fF
C1 sky130_fd_sc_hvl__schmittbuf_1_0/X VSUBS 0.22fF
C2 sky130_fd_sc_hvl__schmittbuf_1_0/A VSUBS 0.49fF
C3 sky130_fd_sc_hvl__schmittbuf_1_0/VPWR VSUBS 0.40fF
C4 sky130_fd_sc_hvl__schmittbuf_1_0/VPB VSUBS 2.88fF
C5 sky130_fd_sc_hvl__schmittbuf_1_0/a_217_207# VSUBS 0.13fF $ **FLOATING
C6 sky130_fd_sc_hvl__schmittbuf_1_0/a_231_463# VSUBS 0.24fF $ **FLOATING
C7 sky130_fd_sc_hvl__schmittbuf_1_0/a_78_463# VSUBS 0.19fF $ **FLOATING
C8 sky130_fd_sc_hvl__schmittbuf_1_0/a_64_207# VSUBS 0.41fF $ **FLOATING
C9 sky130_fd_sc_hvl__schmittbuf_1_0/a_117_181# VSUBS 0.94fF $ **FLOATING
.end

