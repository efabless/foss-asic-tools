magic
tech sky130A
magscale 1 2
timestamp 1624430562
<< error_p >>
rect -1484 566 1484 600
rect -1514 -566 1514 566
rect -1484 -600 1484 -566
<< nwell >>
rect -1484 -600 1484 600
<< mvpmos >>
rect -1390 -500 -1190 500
rect -1132 -500 -932 500
rect -874 -500 -674 500
rect -616 -500 -416 500
rect -358 -500 -158 500
rect -100 -500 100 500
rect 158 -500 358 500
rect 416 -500 616 500
rect 674 -500 874 500
rect 932 -500 1132 500
rect 1190 -500 1390 500
<< mvpdiff >>
rect -1448 488 -1390 500
rect -1448 -488 -1436 488
rect -1402 -488 -1390 488
rect -1448 -500 -1390 -488
rect -1190 488 -1132 500
rect -1190 -488 -1178 488
rect -1144 -488 -1132 488
rect -1190 -500 -1132 -488
rect -932 488 -874 500
rect -932 -488 -920 488
rect -886 -488 -874 488
rect -932 -500 -874 -488
rect -674 488 -616 500
rect -674 -488 -662 488
rect -628 -488 -616 488
rect -674 -500 -616 -488
rect -416 488 -358 500
rect -416 -488 -404 488
rect -370 -488 -358 488
rect -416 -500 -358 -488
rect -158 488 -100 500
rect -158 -488 -146 488
rect -112 -488 -100 488
rect -158 -500 -100 -488
rect 100 488 158 500
rect 100 -488 112 488
rect 146 -488 158 488
rect 100 -500 158 -488
rect 358 488 416 500
rect 358 -488 370 488
rect 404 -488 416 488
rect 358 -500 416 -488
rect 616 488 674 500
rect 616 -488 628 488
rect 662 -488 674 488
rect 616 -500 674 -488
rect 874 488 932 500
rect 874 -488 886 488
rect 920 -488 932 488
rect 874 -500 932 -488
rect 1132 488 1190 500
rect 1132 -488 1144 488
rect 1178 -488 1190 488
rect 1132 -500 1190 -488
rect 1390 488 1448 500
rect 1390 -488 1402 488
rect 1436 -488 1448 488
rect 1390 -500 1448 -488
<< mvpdiffc >>
rect -1436 -488 -1402 488
rect -1178 -488 -1144 488
rect -920 -488 -886 488
rect -662 -488 -628 488
rect -404 -488 -370 488
rect -146 -488 -112 488
rect 112 -488 146 488
rect 370 -488 404 488
rect 628 -488 662 488
rect 886 -488 920 488
rect 1144 -488 1178 488
rect 1402 -488 1436 488
<< poly >>
rect -1356 581 -1224 597
rect -1356 564 -1340 581
rect -1390 547 -1340 564
rect -1240 564 -1224 581
rect -1098 581 -966 597
rect -1098 564 -1082 581
rect -1240 547 -1190 564
rect -1390 500 -1190 547
rect -1132 547 -1082 564
rect -982 564 -966 581
rect -840 581 -708 597
rect -840 564 -824 581
rect -982 547 -932 564
rect -1132 500 -932 547
rect -874 547 -824 564
rect -724 564 -708 581
rect -582 581 -450 597
rect -582 564 -566 581
rect -724 547 -674 564
rect -874 500 -674 547
rect -616 547 -566 564
rect -466 564 -450 581
rect -324 581 -192 597
rect -324 564 -308 581
rect -466 547 -416 564
rect -616 500 -416 547
rect -358 547 -308 564
rect -208 564 -192 581
rect -66 581 66 597
rect -66 564 -50 581
rect -208 547 -158 564
rect -358 500 -158 547
rect -100 547 -50 564
rect 50 564 66 581
rect 192 581 324 597
rect 192 564 208 581
rect 50 547 100 564
rect -100 500 100 547
rect 158 547 208 564
rect 308 564 324 581
rect 450 581 582 597
rect 450 564 466 581
rect 308 547 358 564
rect 158 500 358 547
rect 416 547 466 564
rect 566 564 582 581
rect 708 581 840 597
rect 708 564 724 581
rect 566 547 616 564
rect 416 500 616 547
rect 674 547 724 564
rect 824 564 840 581
rect 966 581 1098 597
rect 966 564 982 581
rect 824 547 874 564
rect 674 500 874 547
rect 932 547 982 564
rect 1082 564 1098 581
rect 1224 581 1356 597
rect 1224 564 1240 581
rect 1082 547 1132 564
rect 932 500 1132 547
rect 1190 547 1240 564
rect 1340 564 1356 581
rect 1340 547 1390 564
rect 1190 500 1390 547
rect -1390 -547 -1190 -500
rect -1390 -564 -1340 -547
rect -1356 -581 -1340 -564
rect -1240 -564 -1190 -547
rect -1132 -547 -932 -500
rect -1132 -564 -1082 -547
rect -1240 -581 -1224 -564
rect -1356 -597 -1224 -581
rect -1098 -581 -1082 -564
rect -982 -564 -932 -547
rect -874 -547 -674 -500
rect -874 -564 -824 -547
rect -982 -581 -966 -564
rect -1098 -597 -966 -581
rect -840 -581 -824 -564
rect -724 -564 -674 -547
rect -616 -547 -416 -500
rect -616 -564 -566 -547
rect -724 -581 -708 -564
rect -840 -597 -708 -581
rect -582 -581 -566 -564
rect -466 -564 -416 -547
rect -358 -547 -158 -500
rect -358 -564 -308 -547
rect -466 -581 -450 -564
rect -582 -597 -450 -581
rect -324 -581 -308 -564
rect -208 -564 -158 -547
rect -100 -547 100 -500
rect -100 -564 -50 -547
rect -208 -581 -192 -564
rect -324 -597 -192 -581
rect -66 -581 -50 -564
rect 50 -564 100 -547
rect 158 -547 358 -500
rect 158 -564 208 -547
rect 50 -581 66 -564
rect -66 -597 66 -581
rect 192 -581 208 -564
rect 308 -564 358 -547
rect 416 -547 616 -500
rect 416 -564 466 -547
rect 308 -581 324 -564
rect 192 -597 324 -581
rect 450 -581 466 -564
rect 566 -564 616 -547
rect 674 -547 874 -500
rect 674 -564 724 -547
rect 566 -581 582 -564
rect 450 -597 582 -581
rect 708 -581 724 -564
rect 824 -564 874 -547
rect 932 -547 1132 -500
rect 932 -564 982 -547
rect 824 -581 840 -564
rect 708 -597 840 -581
rect 966 -581 982 -564
rect 1082 -564 1132 -547
rect 1190 -547 1390 -500
rect 1190 -564 1240 -547
rect 1082 -581 1098 -564
rect 966 -597 1098 -581
rect 1224 -581 1240 -564
rect 1340 -564 1390 -547
rect 1340 -581 1356 -564
rect 1224 -597 1356 -581
<< polycont >>
rect -1340 547 -1240 581
rect -1082 547 -982 581
rect -824 547 -724 581
rect -566 547 -466 581
rect -308 547 -208 581
rect -50 547 50 581
rect 208 547 308 581
rect 466 547 566 581
rect 724 547 824 581
rect 982 547 1082 581
rect 1240 547 1340 581
rect -1340 -581 -1240 -547
rect -1082 -581 -982 -547
rect -824 -581 -724 -547
rect -566 -581 -466 -547
rect -308 -581 -208 -547
rect -50 -581 50 -547
rect 208 -581 308 -547
rect 466 -581 566 -547
rect 724 -581 824 -547
rect 982 -581 1082 -547
rect 1240 -581 1340 -547
<< locali >>
rect -1356 547 -1340 581
rect -1240 547 -1224 581
rect -1098 547 -1082 581
rect -982 547 -966 581
rect -840 547 -824 581
rect -724 547 -708 581
rect -582 547 -566 581
rect -466 547 -450 581
rect -324 547 -308 581
rect -208 547 -192 581
rect -66 547 -50 581
rect 50 547 66 581
rect 192 547 208 581
rect 308 547 324 581
rect 450 547 466 581
rect 566 547 582 581
rect 708 547 724 581
rect 824 547 840 581
rect 966 547 982 581
rect 1082 547 1098 581
rect 1224 547 1240 581
rect 1340 547 1356 581
rect -1436 488 -1402 504
rect -1436 -504 -1402 -488
rect -1178 488 -1144 504
rect -1178 -504 -1144 -488
rect -920 488 -886 504
rect -920 -504 -886 -488
rect -662 488 -628 504
rect -662 -504 -628 -488
rect -404 488 -370 504
rect -404 -504 -370 -488
rect -146 488 -112 504
rect -146 -504 -112 -488
rect 112 488 146 504
rect 112 -504 146 -488
rect 370 488 404 504
rect 370 -504 404 -488
rect 628 488 662 504
rect 628 -504 662 -488
rect 886 488 920 504
rect 886 -504 920 -488
rect 1144 488 1178 504
rect 1144 -504 1178 -488
rect 1402 488 1436 504
rect 1402 -504 1436 -488
rect -1356 -581 -1340 -547
rect -1240 -581 -1224 -547
rect -1098 -581 -1082 -547
rect -982 -581 -966 -547
rect -840 -581 -824 -547
rect -724 -581 -708 -547
rect -582 -581 -566 -547
rect -466 -581 -450 -547
rect -324 -581 -308 -547
rect -208 -581 -192 -547
rect -66 -581 -50 -547
rect 50 -581 66 -547
rect 192 -581 208 -547
rect 308 -581 324 -547
rect 450 -581 466 -547
rect 566 -581 582 -547
rect 708 -581 724 -547
rect 824 -581 840 -547
rect 966 -581 982 -547
rect 1082 -581 1098 -547
rect 1224 -581 1240 -547
rect 1340 -581 1356 -547
<< viali >>
rect -1324 547 -1256 581
rect -1066 547 -998 581
rect -808 547 -740 581
rect -550 547 -482 581
rect -292 547 -224 581
rect -34 547 34 581
rect 224 547 292 581
rect 482 547 550 581
rect 740 547 808 581
rect 998 547 1066 581
rect 1256 547 1324 581
rect -1436 -488 -1402 488
rect -1178 -488 -1144 488
rect -920 -488 -886 488
rect -662 -488 -628 488
rect -404 -488 -370 488
rect -146 -488 -112 488
rect 112 -488 146 488
rect 370 -488 404 488
rect 628 -488 662 488
rect 886 -488 920 488
rect 1144 -488 1178 488
rect 1402 -488 1436 488
rect -1324 -581 -1256 -547
rect -1066 -581 -998 -547
rect -808 -581 -740 -547
rect -550 -581 -482 -547
rect -292 -581 -224 -547
rect -34 -581 34 -547
rect 224 -581 292 -547
rect 482 -581 550 -547
rect 740 -581 808 -547
rect 998 -581 1066 -547
rect 1256 -581 1324 -547
<< metal1 >>
rect -1336 581 -1244 587
rect -1336 547 -1324 581
rect -1256 547 -1244 581
rect -1336 541 -1244 547
rect -1078 581 -986 587
rect -1078 547 -1066 581
rect -998 547 -986 581
rect -1078 541 -986 547
rect -820 581 -728 587
rect -820 547 -808 581
rect -740 547 -728 581
rect -820 541 -728 547
rect -562 581 -470 587
rect -562 547 -550 581
rect -482 547 -470 581
rect -562 541 -470 547
rect -304 581 -212 587
rect -304 547 -292 581
rect -224 547 -212 581
rect -304 541 -212 547
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect 212 581 304 587
rect 212 547 224 581
rect 292 547 304 581
rect 212 541 304 547
rect 470 581 562 587
rect 470 547 482 581
rect 550 547 562 581
rect 470 541 562 547
rect 728 581 820 587
rect 728 547 740 581
rect 808 547 820 581
rect 728 541 820 547
rect 986 581 1078 587
rect 986 547 998 581
rect 1066 547 1078 581
rect 986 541 1078 547
rect 1244 581 1336 587
rect 1244 547 1256 581
rect 1324 547 1336 581
rect 1244 541 1336 547
rect -1442 488 -1396 500
rect -1442 -488 -1436 488
rect -1402 -488 -1396 488
rect -1442 -500 -1396 -488
rect -1184 488 -1138 500
rect -1184 -488 -1178 488
rect -1144 -488 -1138 488
rect -1184 -500 -1138 -488
rect -926 488 -880 500
rect -926 -488 -920 488
rect -886 -488 -880 488
rect -926 -500 -880 -488
rect -668 488 -622 500
rect -668 -488 -662 488
rect -628 -488 -622 488
rect -668 -500 -622 -488
rect -410 488 -364 500
rect -410 -488 -404 488
rect -370 -488 -364 488
rect -410 -500 -364 -488
rect -152 488 -106 500
rect -152 -488 -146 488
rect -112 -488 -106 488
rect -152 -500 -106 -488
rect 106 488 152 500
rect 106 -488 112 488
rect 146 -488 152 488
rect 106 -500 152 -488
rect 364 488 410 500
rect 364 -488 370 488
rect 404 -488 410 488
rect 364 -500 410 -488
rect 622 488 668 500
rect 622 -488 628 488
rect 662 -488 668 488
rect 622 -500 668 -488
rect 880 488 926 500
rect 880 -488 886 488
rect 920 -488 926 488
rect 880 -500 926 -488
rect 1138 488 1184 500
rect 1138 -488 1144 488
rect 1178 -488 1184 488
rect 1138 -500 1184 -488
rect 1396 488 1442 500
rect 1396 -488 1402 488
rect 1436 -488 1442 488
rect 1396 -500 1442 -488
rect -1336 -547 -1244 -541
rect -1336 -581 -1324 -547
rect -1256 -581 -1244 -547
rect -1336 -587 -1244 -581
rect -1078 -547 -986 -541
rect -1078 -581 -1066 -547
rect -998 -581 -986 -547
rect -1078 -587 -986 -581
rect -820 -547 -728 -541
rect -820 -581 -808 -547
rect -740 -581 -728 -547
rect -820 -587 -728 -581
rect -562 -547 -470 -541
rect -562 -581 -550 -547
rect -482 -581 -470 -547
rect -562 -587 -470 -581
rect -304 -547 -212 -541
rect -304 -581 -292 -547
rect -224 -581 -212 -547
rect -304 -587 -212 -581
rect -46 -547 46 -541
rect -46 -581 -34 -547
rect 34 -581 46 -547
rect -46 -587 46 -581
rect 212 -547 304 -541
rect 212 -581 224 -547
rect 292 -581 304 -547
rect 212 -587 304 -581
rect 470 -547 562 -541
rect 470 -581 482 -547
rect 550 -581 562 -547
rect 470 -587 562 -581
rect 728 -547 820 -541
rect 728 -581 740 -547
rect 808 -581 820 -547
rect 728 -587 820 -581
rect 986 -547 1078 -541
rect 986 -581 998 -547
rect 1066 -581 1078 -547
rect 986 -587 1078 -581
rect 1244 -547 1336 -541
rect 1244 -581 1256 -547
rect 1324 -581 1336 -547
rect 1244 -587 1336 -581
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 5 l 1 m 1 nf 11 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
