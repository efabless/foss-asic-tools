magic
tech sky130A
magscale 1 2
timestamp 1624430562
<< nwell >>
rect -8500 0 7600 4000
<< pwell >>
rect -8500 -2400 7600 0
<< mvpsubdiff >>
rect -8400 -124 7500 -100
rect -8400 -2276 -8376 -124
rect -8324 -200 7424 -176
rect -8324 -2200 -8300 -200
rect 7400 -2200 7424 -200
rect -8324 -2224 7424 -2200
rect 7476 -2276 7500 -124
rect -8400 -2300 7500 -2276
<< mvnsubdiff >>
rect -8400 3876 7500 3900
rect -8400 124 -8376 3876
rect -8324 3800 7424 3824
rect -8324 200 -8300 3800
rect 7400 200 7424 3800
rect -8324 176 7424 200
rect 7476 124 7500 3876
rect -8400 100 7500 124
<< mvpsubdiffcont >>
rect -8376 -176 7476 -124
rect -8376 -2224 -8324 -176
rect 7424 -2224 7476 -176
rect -8376 -2276 7476 -2224
<< mvnsubdiffcont >>
rect -8376 3824 7476 3876
rect -8376 176 -8324 3824
rect 7424 176 7476 3824
rect -8376 124 7476 176
<< locali >>
rect -8400 3876 7500 3900
rect -8400 124 -8376 3876
rect -8324 3800 7424 3824
rect -8324 200 -8300 3800
rect -7839 410 -7581 417
rect -7839 370 -7641 410
rect -7595 370 -7581 410
rect -7839 364 -7581 370
rect -7529 364 -7265 417
rect -7529 326 -7423 364
rect -7529 285 -7517 326
rect -7464 285 -7423 326
rect -7529 279 -7423 285
rect 7400 200 7424 3800
rect -8324 191 7424 200
rect -8324 176 -7247 191
rect -6943 188 7424 191
rect -6943 176 -6021 188
rect -5987 176 -4757 188
rect -4723 176 -3493 188
rect -3459 184 -1281 188
rect -3459 176 -2545 184
rect -2511 176 -1281 184
rect -1247 176 -17 188
rect 17 176 1247 188
rect 1281 176 2511 188
rect 2545 176 3775 188
rect 3809 176 5039 188
rect 5073 176 6303 188
rect 6337 176 7424 188
rect 7476 124 7500 3876
rect -8400 100 7500 124
rect -8400 -124 7500 -100
rect -8400 -2276 -8376 -124
rect -8324 -189 -7237 -176
rect -6949 -189 -6021 -176
rect -8324 -190 -6021 -189
rect -5987 -190 -4757 -176
rect -4723 -190 -3493 -176
rect -3459 -190 -2545 -176
rect -2511 -190 -1281 -176
rect -1247 -190 -17 -176
rect 17 -190 1247 -176
rect 1281 -190 2511 -176
rect 2545 -190 3775 -176
rect 3809 -190 5039 -176
rect 5073 -190 6303 -176
rect 6337 -190 7424 -176
rect -8324 -200 7424 -190
rect -8324 -2200 -8300 -200
rect -7789 -901 -7631 -893
rect -7789 -943 -7739 -901
rect -7681 -943 -7631 -901
rect -7789 -974 -7631 -943
rect -7473 -901 -7315 -893
rect -7473 -943 -7423 -901
rect -7366 -943 -7315 -901
rect -7473 -974 -7315 -943
rect 7400 -2200 7424 -200
rect -8324 -2224 7424 -2200
rect 7476 -2276 7500 -124
rect -8400 -2300 7500 -2276
<< viali >>
rect -8376 3824 7476 3876
rect -8376 124 -8324 3824
rect -6890 3511 -6856 3545
rect -6732 3511 -6698 3545
rect -6574 3511 -6540 3545
rect -6416 3511 -6382 3545
rect -6258 3511 -6224 3545
rect -6100 3511 -6066 3545
rect -5942 3511 -5908 3545
rect -5784 3511 -5750 3545
rect -5626 3511 -5592 3545
rect -5468 3511 -5434 3545
rect -5310 3511 -5276 3545
rect -5152 3511 -5118 3545
rect -4994 3511 -4960 3545
rect -4836 3511 -4802 3545
rect -4678 3511 -4644 3545
rect -4520 3511 -4486 3545
rect -4362 3511 -4328 3545
rect -4204 3511 -4170 3545
rect -4046 3511 -4012 3545
rect -3888 3511 -3854 3545
rect -3730 3511 -3696 3545
rect -3572 3511 -3538 3545
rect -3414 3511 -3380 3545
rect -3256 3511 -3222 3545
rect -3098 3511 -3064 3545
rect -2940 3511 -2906 3545
rect -2782 3511 -2748 3545
rect -2624 3511 -2590 3545
rect -2466 3511 -2432 3545
rect -2308 3511 -2274 3545
rect -2150 3511 -2116 3545
rect -1992 3511 -1958 3545
rect -1834 3511 -1800 3545
rect -1676 3511 -1642 3545
rect -1518 3511 -1484 3545
rect -1360 3511 -1326 3545
rect -1202 3511 -1168 3545
rect -1044 3511 -1010 3545
rect -886 3511 -852 3545
rect -728 3511 -694 3545
rect -570 3511 -536 3545
rect -412 3511 -378 3545
rect -254 3511 -220 3545
rect -96 3511 -62 3545
rect 62 3511 96 3545
rect 220 3511 254 3545
rect 378 3511 412 3545
rect 536 3511 570 3545
rect 694 3511 728 3545
rect 852 3511 886 3545
rect 1010 3511 1044 3545
rect 1168 3511 1202 3545
rect 1326 3511 1360 3545
rect 1484 3511 1518 3545
rect 1642 3511 1676 3545
rect 1800 3511 1834 3545
rect 1958 3511 1992 3545
rect 2116 3511 2150 3545
rect 2274 3511 2308 3545
rect 2432 3511 2466 3545
rect 2590 3511 2624 3545
rect 2748 3511 2782 3545
rect 2906 3511 2940 3545
rect 3064 3511 3098 3545
rect 3222 3511 3256 3545
rect 3380 3511 3414 3545
rect 3538 3511 3572 3545
rect 3696 3511 3730 3545
rect 3854 3511 3888 3545
rect 4012 3511 4046 3545
rect 4170 3511 4204 3545
rect 4328 3511 4362 3545
rect 4486 3511 4520 3545
rect 4644 3511 4678 3545
rect 4802 3511 4836 3545
rect 4960 3511 4994 3545
rect 5118 3511 5152 3545
rect 5276 3511 5310 3545
rect 5434 3511 5468 3545
rect 5592 3511 5626 3545
rect 5750 3511 5784 3545
rect 5908 3511 5942 3545
rect 6066 3511 6100 3545
rect 6224 3511 6258 3545
rect 6382 3511 6416 3545
rect 6540 3511 6574 3545
rect 6698 3511 6732 3545
rect 6856 3511 6890 3545
rect -7641 370 -7595 410
rect -6890 383 -6856 417
rect -6732 383 -6698 417
rect -6574 383 -6540 417
rect -6416 383 -6382 417
rect -6258 383 -6224 417
rect -6100 383 -6066 417
rect -5942 383 -5908 417
rect -5784 383 -5750 417
rect -5626 383 -5592 417
rect -5468 383 -5434 417
rect -5310 383 -5276 417
rect -5152 383 -5118 417
rect -4994 383 -4960 417
rect -4836 383 -4802 417
rect -4678 383 -4644 417
rect -4520 383 -4486 417
rect -4362 383 -4328 417
rect -4204 383 -4170 417
rect -4046 383 -4012 417
rect -3888 383 -3854 417
rect -3730 383 -3696 417
rect -3572 383 -3538 417
rect -3414 383 -3380 417
rect -3256 383 -3222 417
rect -3098 383 -3064 417
rect -2940 383 -2906 417
rect -2782 383 -2748 417
rect -2624 383 -2590 417
rect -2466 383 -2432 417
rect -2308 383 -2274 417
rect -2150 383 -2116 417
rect -1992 383 -1958 417
rect -1834 383 -1800 417
rect -1676 383 -1642 417
rect -1518 383 -1484 417
rect -1360 383 -1326 417
rect -1202 383 -1168 417
rect -1044 383 -1010 417
rect -886 383 -852 417
rect -728 383 -694 417
rect -570 383 -536 417
rect -412 383 -378 417
rect -254 383 -220 417
rect -96 383 -62 417
rect 62 383 96 417
rect 220 383 254 417
rect 378 383 412 417
rect 536 383 570 417
rect 694 383 728 417
rect 852 383 886 417
rect 1010 383 1044 417
rect 1168 383 1202 417
rect 1326 383 1360 417
rect 1484 383 1518 417
rect 1642 383 1676 417
rect 1800 383 1834 417
rect 1958 383 1992 417
rect 2116 383 2150 417
rect 2274 383 2308 417
rect 2432 383 2466 417
rect 2590 383 2624 417
rect 2748 383 2782 417
rect 2906 383 2940 417
rect 3064 383 3098 417
rect 3222 383 3256 417
rect 3380 383 3414 417
rect 3538 383 3572 417
rect 3696 383 3730 417
rect 3854 383 3888 417
rect 4012 383 4046 417
rect 4170 383 4204 417
rect 4328 383 4362 417
rect 4486 383 4520 417
rect 4644 383 4678 417
rect 4802 383 4836 417
rect 4960 383 4994 417
rect 5118 383 5152 417
rect 5276 383 5310 417
rect 5434 383 5468 417
rect 5592 383 5626 417
rect 5750 383 5784 417
rect 5908 383 5942 417
rect 6066 383 6100 417
rect 6224 383 6258 417
rect 6382 383 6416 417
rect 6540 383 6574 417
rect 6698 383 6732 417
rect 6856 383 6890 417
rect -7517 285 -7464 326
rect -7247 176 -6943 191
rect -6021 176 -5987 188
rect -4757 176 -4723 188
rect -3493 176 -3459 188
rect -2545 176 -2511 184
rect -1281 176 -1247 188
rect -17 176 17 188
rect 1247 176 1281 188
rect 2511 176 2545 188
rect 3775 176 3809 188
rect 5039 176 5073 188
rect 6303 176 6337 188
rect -7247 145 -6943 176
rect -6021 151 -5987 176
rect -4757 151 -4723 176
rect -3493 151 -3459 176
rect -2545 136 -2511 176
rect -1281 151 -1247 176
rect -17 151 17 176
rect 1247 151 1281 176
rect 2511 151 2545 176
rect 3775 151 3809 176
rect 5039 151 5073 176
rect 6303 151 6337 176
rect 7424 124 7476 3824
rect -8376 -2224 -8324 -124
rect -7237 -176 -6949 -151
rect -6021 -176 -5987 -152
rect -4757 -176 -4723 -152
rect -3493 -176 -3459 -152
rect -2545 -176 -2511 -152
rect -1281 -176 -1247 -152
rect -17 -176 17 -152
rect 1247 -176 1281 -152
rect 2511 -176 2545 -152
rect 3775 -176 3809 -152
rect 5039 -176 5073 -152
rect 6303 -176 6337 -152
rect -7237 -189 -6949 -176
rect -6021 -190 -5987 -176
rect -4757 -190 -4723 -176
rect -3493 -190 -3459 -176
rect -2545 -190 -2511 -176
rect -1281 -190 -1247 -176
rect -17 -190 17 -176
rect 1247 -190 1281 -176
rect 2511 -190 2545 -176
rect 3775 -190 3809 -176
rect 5039 -190 5073 -176
rect 6303 -190 6337 -176
rect -6890 -417 -6856 -383
rect -6732 -417 -6698 -383
rect -6574 -417 -6540 -383
rect -6416 -417 -6382 -383
rect -6258 -417 -6224 -383
rect -6100 -417 -6066 -383
rect -5942 -417 -5908 -383
rect -5784 -417 -5750 -383
rect -5626 -417 -5592 -383
rect -5468 -417 -5434 -383
rect -5310 -417 -5276 -383
rect -5152 -417 -5118 -383
rect -4994 -417 -4960 -383
rect -4836 -417 -4802 -383
rect -4678 -417 -4644 -383
rect -4520 -417 -4486 -383
rect -4362 -417 -4328 -383
rect -4204 -417 -4170 -383
rect -4046 -417 -4012 -383
rect -3888 -417 -3854 -383
rect -3730 -417 -3696 -383
rect -3572 -417 -3538 -383
rect -3414 -417 -3380 -383
rect -3256 -417 -3222 -383
rect -3098 -417 -3064 -383
rect -2940 -417 -2906 -383
rect -2782 -417 -2748 -383
rect -2624 -417 -2590 -383
rect -2466 -417 -2432 -383
rect -2308 -417 -2274 -383
rect -2150 -417 -2116 -383
rect -1992 -417 -1958 -383
rect -1834 -417 -1800 -383
rect -1676 -417 -1642 -383
rect -1518 -417 -1484 -383
rect -1360 -417 -1326 -383
rect -1202 -417 -1168 -383
rect -1044 -417 -1010 -383
rect -886 -417 -852 -383
rect -728 -417 -694 -383
rect -570 -417 -536 -383
rect -412 -417 -378 -383
rect -254 -417 -220 -383
rect -96 -417 -62 -383
rect 62 -417 96 -383
rect 220 -417 254 -383
rect 378 -417 412 -383
rect 536 -417 570 -383
rect 694 -417 728 -383
rect 852 -417 886 -383
rect 1010 -417 1044 -383
rect 1168 -417 1202 -383
rect 1326 -417 1360 -383
rect 1484 -417 1518 -383
rect 1642 -417 1676 -383
rect 1800 -417 1834 -383
rect 1958 -417 1992 -383
rect 2116 -417 2150 -383
rect 2274 -417 2308 -383
rect 2432 -417 2466 -383
rect 2590 -417 2624 -383
rect 2748 -417 2782 -383
rect 2906 -417 2940 -383
rect 3064 -417 3098 -383
rect 3222 -417 3256 -383
rect 3380 -417 3414 -383
rect 3538 -417 3572 -383
rect 3696 -417 3730 -383
rect 3854 -417 3888 -383
rect 4012 -417 4046 -383
rect 4170 -417 4204 -383
rect 4328 -417 4362 -383
rect 4486 -417 4520 -383
rect 4644 -417 4678 -383
rect 4802 -417 4836 -383
rect 4960 -417 4994 -383
rect 5118 -417 5152 -383
rect 5276 -417 5310 -383
rect 5434 -417 5468 -383
rect 5592 -417 5626 -383
rect 5750 -417 5784 -383
rect 5908 -417 5942 -383
rect 6066 -417 6100 -383
rect 6224 -417 6258 -383
rect 6382 -417 6416 -383
rect 6540 -417 6574 -383
rect 6698 -417 6732 -383
rect 6856 -417 6890 -383
rect -7739 -943 -7681 -901
rect -7423 -943 -7366 -901
rect -6890 -1927 -6856 -1893
rect -6732 -1927 -6698 -1893
rect -6574 -1927 -6540 -1893
rect -6416 -1927 -6382 -1893
rect -6258 -1927 -6224 -1893
rect -6100 -1927 -6066 -1893
rect -5942 -1927 -5908 -1893
rect -5784 -1927 -5750 -1893
rect -5626 -1927 -5592 -1893
rect -5468 -1927 -5434 -1893
rect -5310 -1927 -5276 -1893
rect -5152 -1927 -5118 -1893
rect -4994 -1927 -4960 -1893
rect -4836 -1927 -4802 -1893
rect -4678 -1927 -4644 -1893
rect -4520 -1927 -4486 -1893
rect -4362 -1927 -4328 -1893
rect -4204 -1927 -4170 -1893
rect -4046 -1927 -4012 -1893
rect -3888 -1927 -3854 -1893
rect -3730 -1927 -3696 -1893
rect -3572 -1927 -3538 -1893
rect -3414 -1927 -3380 -1893
rect -3256 -1927 -3222 -1893
rect -3098 -1927 -3064 -1893
rect -2940 -1927 -2906 -1893
rect -2782 -1927 -2748 -1893
rect -2624 -1927 -2590 -1893
rect -2466 -1927 -2432 -1893
rect -2308 -1927 -2274 -1893
rect -2150 -1927 -2116 -1893
rect -1992 -1927 -1958 -1893
rect -1834 -1927 -1800 -1893
rect -1676 -1927 -1642 -1893
rect -1518 -1927 -1484 -1893
rect -1360 -1927 -1326 -1893
rect -1202 -1927 -1168 -1893
rect -1044 -1927 -1010 -1893
rect -886 -1927 -852 -1893
rect -728 -1927 -694 -1893
rect -570 -1927 -536 -1893
rect -412 -1927 -378 -1893
rect -254 -1927 -220 -1893
rect -96 -1927 -62 -1893
rect 62 -1927 96 -1893
rect 220 -1927 254 -1893
rect 378 -1927 412 -1893
rect 536 -1927 570 -1893
rect 694 -1927 728 -1893
rect 852 -1927 886 -1893
rect 1010 -1927 1044 -1893
rect 1168 -1927 1202 -1893
rect 1326 -1927 1360 -1893
rect 1484 -1927 1518 -1893
rect 1642 -1927 1676 -1893
rect 1800 -1927 1834 -1893
rect 1958 -1927 1992 -1893
rect 2116 -1927 2150 -1893
rect 2274 -1927 2308 -1893
rect 2432 -1927 2466 -1893
rect 2590 -1927 2624 -1893
rect 2748 -1927 2782 -1893
rect 2906 -1927 2940 -1893
rect 3064 -1927 3098 -1893
rect 3222 -1927 3256 -1893
rect 3380 -1927 3414 -1893
rect 3538 -1927 3572 -1893
rect 3696 -1927 3730 -1893
rect 3854 -1927 3888 -1893
rect 4012 -1927 4046 -1893
rect 4170 -1927 4204 -1893
rect 4328 -1927 4362 -1893
rect 4486 -1927 4520 -1893
rect 4644 -1927 4678 -1893
rect 4802 -1927 4836 -1893
rect 4960 -1927 4994 -1893
rect 5118 -1927 5152 -1893
rect 5276 -1927 5310 -1893
rect 5434 -1927 5468 -1893
rect 5592 -1927 5626 -1893
rect 5750 -1927 5784 -1893
rect 5908 -1927 5942 -1893
rect 6066 -1927 6100 -1893
rect 6224 -1927 6258 -1893
rect 6382 -1927 6416 -1893
rect 6540 -1927 6574 -1893
rect 6698 -1927 6732 -1893
rect 6856 -1927 6890 -1893
rect 7424 -2224 7476 -124
rect -8376 -2276 7476 -2224
<< metal1 >>
rect -8500 3876 7600 4000
rect -8500 3600 -8376 3876
rect -8400 124 -8376 3600
rect -8324 3600 7424 3824
rect -8324 124 -8300 3600
rect -7891 1426 -7213 3600
rect -6975 3464 -6929 3600
rect -6896 3545 -6850 3557
rect -6896 3511 -6890 3545
rect -6856 3511 -6850 3545
rect -7891 1264 -7845 1426
rect -7575 1264 -7529 1426
rect -7259 1264 -7213 1426
rect -8400 100 -8300 124
rect -7733 336 -7687 464
rect -7417 417 -7371 464
rect -7653 410 -7371 417
rect -7653 370 -7641 410
rect -7595 370 -7371 410
rect -7653 364 -7371 370
rect -7733 326 -7451 336
rect -7733 285 -7517 326
rect -7464 285 -7451 326
rect -7733 279 -7451 285
rect -8400 -124 -8300 -100
rect -8400 -2000 -8376 -124
rect -8500 -2276 -8376 -2000
rect -8324 -2000 -8300 -124
rect -7733 -455 -7687 279
rect -7417 100 -7371 364
rect -7259 191 -6929 464
rect -7259 145 -7247 191
rect -6943 145 -6929 191
rect -7259 139 -6929 145
rect -6896 417 -6850 3511
rect -6738 3545 -6692 3557
rect -6738 3511 -6732 3545
rect -6698 3511 -6692 3545
rect -6817 446 -6771 464
rect -6896 383 -6890 417
rect -6856 383 -6850 417
rect -6896 100 -6850 383
rect -6820 440 -6768 446
rect -6820 382 -6768 388
rect -6738 417 -6692 3511
rect -6659 3464 -6613 3600
rect -6580 3545 -6534 3557
rect -6580 3511 -6574 3545
rect -6540 3511 -6534 3545
rect -6738 383 -6732 417
rect -6698 383 -6692 417
rect -6738 100 -6692 383
rect -7417 -100 -6692 100
rect -7417 -455 -7371 -100
rect -7259 -151 -6929 -140
rect -7259 -189 -7237 -151
rect -6949 -189 -6929 -151
rect -7259 -455 -6929 -189
rect -6896 -383 -6850 -100
rect -6896 -417 -6890 -383
rect -6856 -417 -6850 -383
rect -7891 -1144 -7845 -855
rect -7789 -901 -7631 -893
rect -7789 -959 -7739 -901
rect -7681 -943 -7631 -901
rect -7682 -959 -7631 -943
rect -7789 -974 -7631 -959
rect -7575 -1144 -7529 -855
rect -7473 -901 -7315 -893
rect -7473 -959 -7423 -901
rect -7366 -959 -7315 -901
rect -7473 -974 -7315 -959
rect -7259 -1144 -7213 -855
rect -7891 -2000 -7213 -1144
rect -6975 -2000 -6929 -1855
rect -6896 -1893 -6850 -417
rect -6820 -379 -6768 -373
rect -6820 -437 -6768 -431
rect -6738 -383 -6692 -100
rect -6738 -417 -6732 -383
rect -6698 -417 -6692 -383
rect -6817 -455 -6771 -437
rect -6896 -1927 -6890 -1893
rect -6856 -1927 -6850 -1893
rect -6896 -1939 -6850 -1927
rect -6738 -1893 -6692 -417
rect -6580 417 -6534 3511
rect -6422 3545 -6376 3557
rect -6422 3511 -6416 3545
rect -6382 3511 -6376 3545
rect -6501 446 -6455 464
rect -6580 383 -6574 417
rect -6540 383 -6534 417
rect -6580 100 -6534 383
rect -6504 440 -6452 446
rect -6504 382 -6452 388
rect -6422 417 -6376 3511
rect -6343 3464 -6297 3600
rect -6264 3545 -6218 3557
rect -6264 3511 -6258 3545
rect -6224 3511 -6218 3545
rect -6422 383 -6416 417
rect -6382 383 -6376 417
rect -6422 100 -6376 383
rect -6264 417 -6218 3511
rect -6106 3545 -6060 3557
rect -6106 3511 -6100 3545
rect -6066 3511 -6060 3545
rect -6185 446 -6139 464
rect -6264 383 -6258 417
rect -6224 383 -6218 417
rect -6264 100 -6218 383
rect -6188 440 -6136 446
rect -6188 382 -6136 388
rect -6106 417 -6060 3511
rect -6027 3464 -5981 3600
rect -5948 3545 -5902 3557
rect -5948 3511 -5942 3545
rect -5908 3511 -5902 3545
rect -6106 383 -6100 417
rect -6066 383 -6060 417
rect -6106 100 -6060 383
rect -6027 188 -5981 464
rect -6027 151 -6021 188
rect -5987 151 -5981 188
rect -6027 139 -5981 151
rect -5948 417 -5902 3511
rect -5790 3545 -5744 3557
rect -5790 3511 -5784 3545
rect -5750 3511 -5744 3545
rect -5869 446 -5823 464
rect -5948 383 -5942 417
rect -5908 383 -5902 417
rect -5948 100 -5902 383
rect -5872 440 -5820 446
rect -5872 382 -5820 388
rect -5790 417 -5744 3511
rect -5711 3464 -5665 3600
rect -5632 3545 -5586 3557
rect -5632 3511 -5626 3545
rect -5592 3511 -5586 3545
rect -5790 383 -5784 417
rect -5750 383 -5744 417
rect -5790 100 -5744 383
rect -6580 80 -5744 100
rect -6580 -80 -6560 80
rect -6246 -80 -5744 80
rect -6580 -100 -5744 -80
rect -6580 -383 -6534 -100
rect -6580 -417 -6574 -383
rect -6540 -417 -6534 -383
rect -6738 -1927 -6732 -1893
rect -6698 -1927 -6692 -1893
rect -6738 -1939 -6692 -1927
rect -6659 -2000 -6613 -1855
rect -6580 -1893 -6534 -417
rect -6504 -379 -6452 -373
rect -6504 -437 -6452 -431
rect -6422 -383 -6376 -100
rect -6422 -417 -6416 -383
rect -6382 -417 -6376 -383
rect -6501 -455 -6455 -437
rect -6580 -1927 -6574 -1893
rect -6540 -1927 -6534 -1893
rect -6580 -1939 -6534 -1927
rect -6422 -1893 -6376 -417
rect -6264 -383 -6218 -100
rect -6264 -417 -6258 -383
rect -6224 -417 -6218 -383
rect -6422 -1927 -6416 -1893
rect -6382 -1927 -6376 -1893
rect -6422 -1939 -6376 -1927
rect -6343 -2000 -6297 -1855
rect -6264 -1893 -6218 -417
rect -6188 -379 -6136 -373
rect -6188 -437 -6136 -431
rect -6106 -383 -6060 -100
rect -6106 -417 -6100 -383
rect -6066 -417 -6060 -383
rect -6185 -455 -6139 -437
rect -6264 -1927 -6258 -1893
rect -6224 -1927 -6218 -1893
rect -6264 -1939 -6218 -1927
rect -6106 -1893 -6060 -417
rect -6027 -152 -5981 -140
rect -6027 -190 -6021 -152
rect -5987 -190 -5981 -152
rect -6027 -455 -5981 -190
rect -5948 -383 -5902 -100
rect -5948 -417 -5942 -383
rect -5908 -417 -5902 -383
rect -6106 -1927 -6100 -1893
rect -6066 -1927 -6060 -1893
rect -6106 -1939 -6060 -1927
rect -6027 -2000 -5981 -1855
rect -5948 -1893 -5902 -417
rect -5872 -379 -5820 -373
rect -5872 -437 -5820 -431
rect -5790 -383 -5744 -100
rect -5790 -417 -5784 -383
rect -5750 -417 -5744 -383
rect -5869 -455 -5823 -437
rect -5948 -1927 -5942 -1893
rect -5908 -1927 -5902 -1893
rect -5948 -1939 -5902 -1927
rect -5790 -1893 -5744 -417
rect -5632 417 -5586 3511
rect -5474 3545 -5428 3557
rect -5474 3511 -5468 3545
rect -5434 3511 -5428 3545
rect -5553 446 -5507 464
rect -5632 383 -5626 417
rect -5592 383 -5586 417
rect -5632 100 -5586 383
rect -5556 440 -5504 446
rect -5556 382 -5504 388
rect -5474 417 -5428 3511
rect -5395 3464 -5349 3600
rect -5316 3545 -5270 3557
rect -5316 3511 -5310 3545
rect -5276 3511 -5270 3545
rect -5474 383 -5468 417
rect -5434 383 -5428 417
rect -5474 100 -5428 383
rect -5316 417 -5270 3511
rect -5158 3545 -5112 3557
rect -5158 3511 -5152 3545
rect -5118 3511 -5112 3545
rect -5237 446 -5191 464
rect -5316 383 -5310 417
rect -5276 383 -5270 417
rect -5316 100 -5270 383
rect -5240 440 -5188 446
rect -5240 382 -5188 388
rect -5158 417 -5112 3511
rect -5079 3464 -5033 3600
rect -5000 3545 -4954 3557
rect -5000 3511 -4994 3545
rect -4960 3511 -4954 3545
rect -5158 383 -5152 417
rect -5118 383 -5112 417
rect -5158 100 -5112 383
rect -5000 417 -4954 3511
rect -4842 3545 -4796 3557
rect -4842 3511 -4836 3545
rect -4802 3511 -4796 3545
rect -4921 446 -4875 464
rect -5000 383 -4994 417
rect -4960 383 -4954 417
rect -5000 100 -4954 383
rect -4924 440 -4872 446
rect -4924 382 -4872 388
rect -4842 417 -4796 3511
rect -4763 3464 -4717 3600
rect -4684 3545 -4638 3557
rect -4684 3511 -4678 3545
rect -4644 3511 -4638 3545
rect -4842 383 -4836 417
rect -4802 383 -4796 417
rect -4842 100 -4796 383
rect -4763 188 -4717 464
rect -4763 151 -4757 188
rect -4723 151 -4717 188
rect -4763 139 -4717 151
rect -4684 417 -4638 3511
rect -4526 3545 -4480 3557
rect -4526 3511 -4520 3545
rect -4486 3511 -4480 3545
rect -4605 446 -4559 464
rect -4684 383 -4678 417
rect -4644 383 -4638 417
rect -4684 100 -4638 383
rect -4608 440 -4556 446
rect -4608 382 -4556 388
rect -4526 417 -4480 3511
rect -4447 3464 -4401 3600
rect -4368 3545 -4322 3557
rect -4368 3511 -4362 3545
rect -4328 3511 -4322 3545
rect -4526 383 -4520 417
rect -4486 383 -4480 417
rect -4526 100 -4480 383
rect -4368 417 -4322 3511
rect -4210 3545 -4164 3557
rect -4210 3511 -4204 3545
rect -4170 3511 -4164 3545
rect -4289 446 -4243 464
rect -4368 383 -4362 417
rect -4328 383 -4322 417
rect -4368 100 -4322 383
rect -4292 440 -4240 446
rect -4292 382 -4240 388
rect -4210 417 -4164 3511
rect -4131 3464 -4085 3600
rect -4052 3545 -4006 3557
rect -4052 3511 -4046 3545
rect -4012 3511 -4006 3545
rect -4210 383 -4204 417
rect -4170 383 -4164 417
rect -4210 100 -4164 383
rect -4052 417 -4006 3511
rect -3894 3545 -3848 3557
rect -3894 3511 -3888 3545
rect -3854 3511 -3848 3545
rect -3973 446 -3927 464
rect -4052 383 -4046 417
rect -4012 383 -4006 417
rect -4052 100 -4006 383
rect -3976 440 -3924 446
rect -3976 382 -3924 388
rect -3894 417 -3848 3511
rect -3815 3464 -3769 3600
rect -3736 3545 -3690 3557
rect -3736 3511 -3730 3545
rect -3696 3511 -3690 3545
rect -3894 383 -3888 417
rect -3854 383 -3848 417
rect -3894 100 -3848 383
rect -3736 417 -3690 3511
rect -3578 3545 -3532 3557
rect -3578 3511 -3572 3545
rect -3538 3511 -3532 3545
rect -3657 446 -3611 464
rect -3736 383 -3730 417
rect -3696 383 -3690 417
rect -3736 100 -3690 383
rect -3660 440 -3608 446
rect -3660 382 -3608 388
rect -3578 417 -3532 3511
rect -3499 3464 -3453 3600
rect -3420 3545 -3374 3557
rect -3420 3511 -3414 3545
rect -3380 3511 -3374 3545
rect -3578 383 -3572 417
rect -3538 383 -3532 417
rect -3578 100 -3532 383
rect -3499 188 -3453 464
rect -3499 151 -3493 188
rect -3459 151 -3453 188
rect -3499 139 -3453 151
rect -3420 417 -3374 3511
rect -3262 3545 -3216 3557
rect -3262 3511 -3256 3545
rect -3222 3511 -3216 3545
rect -3341 446 -3295 464
rect -3420 383 -3414 417
rect -3380 383 -3374 417
rect -3420 100 -3374 383
rect -3344 440 -3292 446
rect -3344 382 -3292 388
rect -3262 417 -3216 3511
rect -3183 3464 -3137 3600
rect -3104 3545 -3058 3557
rect -3104 3511 -3098 3545
rect -3064 3511 -3058 3545
rect -3262 383 -3256 417
rect -3222 383 -3216 417
rect -3262 100 -3216 383
rect -3104 417 -3058 3511
rect -2946 3545 -2900 3557
rect -2946 3511 -2940 3545
rect -2906 3511 -2900 3545
rect -3025 446 -2979 464
rect -3104 383 -3098 417
rect -3064 383 -3058 417
rect -3104 100 -3058 383
rect -3028 440 -2976 446
rect -3028 382 -2976 388
rect -2946 417 -2900 3511
rect -2867 3464 -2821 3600
rect -2788 3545 -2742 3557
rect -2788 3511 -2782 3545
rect -2748 3511 -2742 3545
rect -2946 383 -2940 417
rect -2906 383 -2900 417
rect -2946 100 -2900 383
rect -2788 417 -2742 3511
rect -2630 3545 -2584 3557
rect -2630 3511 -2624 3545
rect -2590 3511 -2584 3545
rect -2709 446 -2663 464
rect -2788 383 -2782 417
rect -2748 383 -2742 417
rect -2788 100 -2742 383
rect -2712 440 -2660 446
rect -2712 382 -2660 388
rect -2630 417 -2584 3511
rect -2551 3464 -2505 3600
rect -2472 3545 -2426 3557
rect -2472 3511 -2466 3545
rect -2432 3511 -2426 3545
rect -2630 383 -2624 417
rect -2590 383 -2584 417
rect -2630 100 -2584 383
rect -2551 184 -2505 464
rect -2551 136 -2545 184
rect -2511 136 -2505 184
rect -2551 124 -2505 136
rect -2472 417 -2426 3511
rect -2314 3545 -2268 3557
rect -2314 3511 -2308 3545
rect -2274 3511 -2268 3545
rect -2393 446 -2347 464
rect -2472 383 -2466 417
rect -2432 383 -2426 417
rect -5632 80 -2584 100
rect -5632 -80 -5562 80
rect -3078 -80 -2584 80
rect -5632 -100 -2584 -80
rect -5632 -383 -5586 -100
rect -5632 -417 -5626 -383
rect -5592 -417 -5586 -383
rect -5790 -1927 -5784 -1893
rect -5750 -1927 -5744 -1893
rect -5790 -1939 -5744 -1927
rect -5711 -2000 -5665 -1855
rect -5632 -1893 -5586 -417
rect -5556 -379 -5504 -373
rect -5556 -437 -5504 -431
rect -5474 -383 -5428 -100
rect -5474 -417 -5468 -383
rect -5434 -417 -5428 -383
rect -5553 -455 -5507 -437
rect -5632 -1927 -5626 -1893
rect -5592 -1927 -5586 -1893
rect -5632 -1939 -5586 -1927
rect -5474 -1893 -5428 -417
rect -5316 -383 -5270 -100
rect -5316 -417 -5310 -383
rect -5276 -417 -5270 -383
rect -5474 -1927 -5468 -1893
rect -5434 -1927 -5428 -1893
rect -5474 -1939 -5428 -1927
rect -5395 -2000 -5349 -1855
rect -5316 -1893 -5270 -417
rect -5240 -379 -5188 -373
rect -5240 -437 -5188 -431
rect -5158 -383 -5112 -100
rect -5158 -417 -5152 -383
rect -5118 -417 -5112 -383
rect -5237 -455 -5191 -437
rect -5316 -1927 -5310 -1893
rect -5276 -1927 -5270 -1893
rect -5316 -1939 -5270 -1927
rect -5158 -1893 -5112 -417
rect -5000 -383 -4954 -100
rect -5000 -417 -4994 -383
rect -4960 -417 -4954 -383
rect -5158 -1927 -5152 -1893
rect -5118 -1927 -5112 -1893
rect -5158 -1939 -5112 -1927
rect -5079 -2000 -5033 -1855
rect -5000 -1893 -4954 -417
rect -4924 -379 -4872 -373
rect -4924 -437 -4872 -431
rect -4842 -383 -4796 -100
rect -4842 -417 -4836 -383
rect -4802 -417 -4796 -383
rect -4921 -455 -4875 -437
rect -5000 -1927 -4994 -1893
rect -4960 -1927 -4954 -1893
rect -5000 -1939 -4954 -1927
rect -4842 -1893 -4796 -417
rect -4763 -152 -4717 -140
rect -4763 -190 -4757 -152
rect -4723 -190 -4717 -152
rect -4763 -455 -4717 -190
rect -4684 -383 -4638 -100
rect -4684 -417 -4678 -383
rect -4644 -417 -4638 -383
rect -4842 -1927 -4836 -1893
rect -4802 -1927 -4796 -1893
rect -4842 -1939 -4796 -1927
rect -4763 -2000 -4717 -1855
rect -4684 -1893 -4638 -417
rect -4608 -379 -4556 -373
rect -4608 -437 -4556 -431
rect -4526 -383 -4480 -100
rect -4526 -417 -4520 -383
rect -4486 -417 -4480 -383
rect -4605 -455 -4559 -437
rect -4684 -1927 -4678 -1893
rect -4644 -1927 -4638 -1893
rect -4684 -1939 -4638 -1927
rect -4526 -1893 -4480 -417
rect -4368 -383 -4322 -100
rect -4368 -417 -4362 -383
rect -4328 -417 -4322 -383
rect -4526 -1927 -4520 -1893
rect -4486 -1927 -4480 -1893
rect -4526 -1939 -4480 -1927
rect -4447 -2000 -4401 -1855
rect -4368 -1893 -4322 -417
rect -4292 -379 -4240 -373
rect -4292 -437 -4240 -431
rect -4210 -383 -4164 -100
rect -4210 -417 -4204 -383
rect -4170 -417 -4164 -383
rect -4289 -455 -4243 -437
rect -4368 -1927 -4362 -1893
rect -4328 -1927 -4322 -1893
rect -4368 -1939 -4322 -1927
rect -4210 -1893 -4164 -417
rect -4052 -383 -4006 -100
rect -4052 -417 -4046 -383
rect -4012 -417 -4006 -383
rect -4210 -1927 -4204 -1893
rect -4170 -1927 -4164 -1893
rect -4210 -1939 -4164 -1927
rect -4131 -2000 -4085 -1855
rect -4052 -1893 -4006 -417
rect -3976 -379 -3924 -373
rect -3976 -437 -3924 -431
rect -3894 -383 -3848 -100
rect -3894 -417 -3888 -383
rect -3854 -417 -3848 -383
rect -3973 -455 -3927 -437
rect -4052 -1927 -4046 -1893
rect -4012 -1927 -4006 -1893
rect -4052 -1939 -4006 -1927
rect -3894 -1893 -3848 -417
rect -3736 -383 -3690 -100
rect -3736 -417 -3730 -383
rect -3696 -417 -3690 -383
rect -3894 -1927 -3888 -1893
rect -3854 -1927 -3848 -1893
rect -3894 -1939 -3848 -1927
rect -3815 -2000 -3769 -1855
rect -3736 -1893 -3690 -417
rect -3660 -379 -3608 -373
rect -3660 -437 -3608 -431
rect -3578 -383 -3532 -100
rect -3578 -417 -3572 -383
rect -3538 -417 -3532 -383
rect -3657 -455 -3611 -437
rect -3736 -1927 -3730 -1893
rect -3696 -1927 -3690 -1893
rect -3736 -1939 -3690 -1927
rect -3578 -1893 -3532 -417
rect -3499 -152 -3453 -140
rect -3499 -190 -3493 -152
rect -3459 -190 -3453 -152
rect -3499 -455 -3453 -190
rect -3420 -383 -3374 -100
rect -3420 -417 -3414 -383
rect -3380 -417 -3374 -383
rect -3578 -1927 -3572 -1893
rect -3538 -1927 -3532 -1893
rect -3578 -1939 -3532 -1927
rect -3499 -2000 -3453 -1855
rect -3420 -1893 -3374 -417
rect -3344 -379 -3292 -373
rect -3344 -437 -3292 -431
rect -3262 -383 -3216 -100
rect -3262 -417 -3256 -383
rect -3222 -417 -3216 -383
rect -3341 -455 -3295 -437
rect -3420 -1927 -3414 -1893
rect -3380 -1927 -3374 -1893
rect -3420 -1939 -3374 -1927
rect -3262 -1893 -3216 -417
rect -3104 -383 -3058 -100
rect -3104 -417 -3098 -383
rect -3064 -417 -3058 -383
rect -3262 -1927 -3256 -1893
rect -3222 -1927 -3216 -1893
rect -3262 -1939 -3216 -1927
rect -3183 -2000 -3137 -1855
rect -3104 -1893 -3058 -417
rect -3028 -379 -2976 -373
rect -3028 -437 -2976 -431
rect -2946 -383 -2900 -100
rect -2946 -417 -2940 -383
rect -2906 -417 -2900 -383
rect -3025 -455 -2979 -437
rect -3104 -1927 -3098 -1893
rect -3064 -1927 -3058 -1893
rect -3104 -1939 -3058 -1927
rect -2946 -1893 -2900 -417
rect -2788 -383 -2742 -100
rect -2788 -417 -2782 -383
rect -2748 -417 -2742 -383
rect -2946 -1927 -2940 -1893
rect -2906 -1927 -2900 -1893
rect -2946 -1939 -2900 -1927
rect -2867 -2000 -2821 -1855
rect -2788 -1893 -2742 -417
rect -2712 -379 -2660 -373
rect -2712 -437 -2660 -431
rect -2630 -383 -2584 -100
rect -2472 100 -2426 383
rect -2396 440 -2344 446
rect -2396 382 -2344 388
rect -2314 417 -2268 3511
rect -2235 3464 -2189 3600
rect -2156 3545 -2110 3557
rect -2156 3511 -2150 3545
rect -2116 3511 -2110 3545
rect -2314 383 -2308 417
rect -2274 383 -2268 417
rect -2314 100 -2268 383
rect -2156 417 -2110 3511
rect -1998 3545 -1952 3557
rect -1998 3511 -1992 3545
rect -1958 3511 -1952 3545
rect -2077 446 -2031 464
rect -2156 383 -2150 417
rect -2116 383 -2110 417
rect -2156 100 -2110 383
rect -2080 440 -2028 446
rect -2080 382 -2028 388
rect -1998 417 -1952 3511
rect -1919 3464 -1873 3600
rect -1840 3545 -1794 3557
rect -1840 3511 -1834 3545
rect -1800 3511 -1794 3545
rect -1998 383 -1992 417
rect -1958 383 -1952 417
rect -1998 100 -1952 383
rect -1840 417 -1794 3511
rect -1682 3545 -1636 3557
rect -1682 3511 -1676 3545
rect -1642 3511 -1636 3545
rect -1761 446 -1715 464
rect -1840 383 -1834 417
rect -1800 383 -1794 417
rect -1840 100 -1794 383
rect -1764 440 -1712 446
rect -1764 382 -1712 388
rect -1682 417 -1636 3511
rect -1603 3464 -1557 3600
rect -1524 3545 -1478 3557
rect -1524 3511 -1518 3545
rect -1484 3511 -1478 3545
rect -1682 383 -1676 417
rect -1642 383 -1636 417
rect -1682 100 -1636 383
rect -1524 417 -1478 3511
rect -1366 3545 -1320 3557
rect -1366 3511 -1360 3545
rect -1326 3511 -1320 3545
rect -1445 446 -1399 464
rect -1524 383 -1518 417
rect -1484 383 -1478 417
rect -1524 100 -1478 383
rect -1448 440 -1396 446
rect -1448 382 -1396 388
rect -1366 417 -1320 3511
rect -1287 3464 -1241 3600
rect -1208 3545 -1162 3557
rect -1208 3511 -1202 3545
rect -1168 3511 -1162 3545
rect -1366 383 -1360 417
rect -1326 383 -1320 417
rect -1366 100 -1320 383
rect -1287 188 -1241 464
rect -1287 151 -1281 188
rect -1247 151 -1241 188
rect -1287 139 -1241 151
rect -1208 417 -1162 3511
rect -1050 3545 -1004 3557
rect -1050 3511 -1044 3545
rect -1010 3511 -1004 3545
rect -1129 446 -1083 464
rect -1208 383 -1202 417
rect -1168 383 -1162 417
rect -1208 100 -1162 383
rect -1132 440 -1080 446
rect -1132 382 -1080 388
rect -1050 417 -1004 3511
rect -971 3464 -925 3600
rect -892 3545 -846 3557
rect -892 3511 -886 3545
rect -852 3511 -846 3545
rect -1050 383 -1044 417
rect -1010 383 -1004 417
rect -1050 100 -1004 383
rect -892 417 -846 3511
rect -734 3545 -688 3557
rect -734 3511 -728 3545
rect -694 3511 -688 3545
rect -813 446 -767 464
rect -892 383 -886 417
rect -852 383 -846 417
rect -892 100 -846 383
rect -816 440 -764 446
rect -816 382 -764 388
rect -734 417 -688 3511
rect -655 3464 -609 3600
rect -576 3545 -530 3557
rect -576 3511 -570 3545
rect -536 3511 -530 3545
rect -734 383 -728 417
rect -694 383 -688 417
rect -734 100 -688 383
rect -576 417 -530 3511
rect -418 3545 -372 3557
rect -418 3511 -412 3545
rect -378 3511 -372 3545
rect -497 446 -451 464
rect -576 383 -570 417
rect -536 383 -530 417
rect -576 100 -530 383
rect -500 440 -448 446
rect -500 382 -448 388
rect -418 417 -372 3511
rect -339 3464 -293 3600
rect -260 3545 -214 3557
rect -260 3511 -254 3545
rect -220 3511 -214 3545
rect -418 383 -412 417
rect -378 383 -372 417
rect -418 100 -372 383
rect -260 417 -214 3511
rect -102 3545 -56 3557
rect -102 3511 -96 3545
rect -62 3511 -56 3545
rect -181 446 -135 464
rect -260 383 -254 417
rect -220 383 -214 417
rect -260 100 -214 383
rect -184 440 -132 446
rect -184 382 -132 388
rect -102 417 -56 3511
rect -23 3464 23 3600
rect 56 3545 102 3557
rect 56 3511 62 3545
rect 96 3511 102 3545
rect -102 383 -96 417
rect -62 383 -56 417
rect -102 100 -56 383
rect -23 188 23 464
rect -23 151 -17 188
rect 17 151 23 188
rect -23 139 23 151
rect 56 417 102 3511
rect 214 3545 260 3557
rect 214 3511 220 3545
rect 254 3511 260 3545
rect 135 446 181 464
rect 56 383 62 417
rect 96 383 102 417
rect 56 100 102 383
rect 132 440 184 446
rect 132 382 184 388
rect 214 417 260 3511
rect 293 3464 339 3600
rect 372 3545 418 3557
rect 372 3511 378 3545
rect 412 3511 418 3545
rect 214 383 220 417
rect 254 383 260 417
rect 214 100 260 383
rect 372 417 418 3511
rect 530 3545 576 3557
rect 530 3511 536 3545
rect 570 3511 576 3545
rect 451 446 497 464
rect 372 383 378 417
rect 412 383 418 417
rect 372 100 418 383
rect 448 440 500 446
rect 448 382 500 388
rect 530 417 576 3511
rect 609 3464 655 3600
rect 688 3545 734 3557
rect 688 3511 694 3545
rect 728 3511 734 3545
rect 530 383 536 417
rect 570 383 576 417
rect 530 100 576 383
rect 688 417 734 3511
rect 846 3545 892 3557
rect 846 3511 852 3545
rect 886 3511 892 3545
rect 767 446 813 464
rect 688 383 694 417
rect 728 383 734 417
rect 688 100 734 383
rect 764 440 816 446
rect 764 382 816 388
rect 846 417 892 3511
rect 925 3464 971 3600
rect 1004 3545 1050 3557
rect 1004 3511 1010 3545
rect 1044 3511 1050 3545
rect 846 383 852 417
rect 886 383 892 417
rect 846 100 892 383
rect 1004 417 1050 3511
rect 1162 3545 1208 3557
rect 1162 3511 1168 3545
rect 1202 3511 1208 3545
rect 1083 446 1129 464
rect 1004 383 1010 417
rect 1044 383 1050 417
rect 1004 100 1050 383
rect 1080 440 1132 446
rect 1080 382 1132 388
rect 1162 417 1208 3511
rect 1241 3464 1287 3600
rect 1320 3545 1366 3557
rect 1320 3511 1326 3545
rect 1360 3511 1366 3545
rect 1162 383 1168 417
rect 1202 383 1208 417
rect 1162 100 1208 383
rect 1241 188 1287 464
rect 1241 151 1247 188
rect 1281 151 1287 188
rect 1241 139 1287 151
rect 1320 417 1366 3511
rect 1478 3545 1524 3557
rect 1478 3511 1484 3545
rect 1518 3511 1524 3545
rect 1399 446 1445 464
rect 1320 383 1326 417
rect 1360 383 1366 417
rect 1320 100 1366 383
rect 1396 440 1448 446
rect 1396 382 1448 388
rect 1478 417 1524 3511
rect 1557 3464 1603 3600
rect 1636 3545 1682 3557
rect 1636 3511 1642 3545
rect 1676 3511 1682 3545
rect 1478 383 1484 417
rect 1518 383 1524 417
rect 1478 100 1524 383
rect 1636 417 1682 3511
rect 1794 3545 1840 3557
rect 1794 3511 1800 3545
rect 1834 3511 1840 3545
rect 1715 446 1761 464
rect 1636 383 1642 417
rect 1676 383 1682 417
rect 1636 100 1682 383
rect 1712 440 1764 446
rect 1712 382 1764 388
rect 1794 417 1840 3511
rect 1873 3464 1919 3600
rect 1952 3545 1998 3557
rect 1952 3511 1958 3545
rect 1992 3511 1998 3545
rect 1794 383 1800 417
rect 1834 383 1840 417
rect 1794 100 1840 383
rect 1952 417 1998 3511
rect 2110 3545 2156 3557
rect 2110 3511 2116 3545
rect 2150 3511 2156 3545
rect 2031 446 2077 464
rect 1952 383 1958 417
rect 1992 383 1998 417
rect 1952 100 1998 383
rect 2028 440 2080 446
rect 2028 382 2080 388
rect 2110 417 2156 3511
rect 2189 3464 2235 3600
rect 2268 3545 2314 3557
rect 2268 3511 2274 3545
rect 2308 3511 2314 3545
rect 2110 383 2116 417
rect 2150 383 2156 417
rect 2110 100 2156 383
rect 2268 417 2314 3511
rect 2426 3545 2472 3557
rect 2426 3511 2432 3545
rect 2466 3511 2472 3545
rect 2347 446 2393 464
rect 2268 383 2274 417
rect 2308 383 2314 417
rect 2268 100 2314 383
rect 2344 440 2396 446
rect 2344 382 2396 388
rect 2426 417 2472 3511
rect 2505 3464 2551 3600
rect 2584 3545 2630 3557
rect 2584 3511 2590 3545
rect 2624 3511 2630 3545
rect 2426 383 2432 417
rect 2466 383 2472 417
rect 2426 100 2472 383
rect 2505 188 2551 464
rect 2505 151 2511 188
rect 2545 151 2551 188
rect 2505 139 2551 151
rect 2584 417 2630 3511
rect 2742 3545 2788 3557
rect 2742 3511 2748 3545
rect 2782 3511 2788 3545
rect 2663 446 2709 464
rect 2584 383 2590 417
rect 2624 383 2630 417
rect 2584 100 2630 383
rect 2660 440 2712 446
rect 2660 382 2712 388
rect 2742 417 2788 3511
rect 2821 3464 2867 3600
rect 2900 3545 2946 3557
rect 2900 3511 2906 3545
rect 2940 3511 2946 3545
rect 2742 383 2748 417
rect 2782 383 2788 417
rect 2742 100 2788 383
rect 2900 417 2946 3511
rect 3058 3545 3104 3557
rect 3058 3511 3064 3545
rect 3098 3511 3104 3545
rect 2979 446 3025 464
rect 2900 383 2906 417
rect 2940 383 2946 417
rect 2900 100 2946 383
rect 2976 440 3028 446
rect 2976 382 3028 388
rect 3058 417 3104 3511
rect 3137 3464 3183 3600
rect 3216 3545 3262 3557
rect 3216 3511 3222 3545
rect 3256 3511 3262 3545
rect 3058 383 3064 417
rect 3098 383 3104 417
rect 3058 100 3104 383
rect 3216 417 3262 3511
rect 3374 3545 3420 3557
rect 3374 3511 3380 3545
rect 3414 3511 3420 3545
rect 3295 446 3341 464
rect 3216 383 3222 417
rect 3256 383 3262 417
rect 3216 100 3262 383
rect 3292 440 3344 446
rect 3292 382 3344 388
rect 3374 417 3420 3511
rect 3453 3464 3499 3600
rect 3532 3545 3578 3557
rect 3532 3511 3538 3545
rect 3572 3511 3578 3545
rect 3374 383 3380 417
rect 3414 383 3420 417
rect 3374 100 3420 383
rect 3532 417 3578 3511
rect 3690 3545 3736 3557
rect 3690 3511 3696 3545
rect 3730 3511 3736 3545
rect 3611 446 3657 464
rect 3532 383 3538 417
rect 3572 383 3578 417
rect 3532 100 3578 383
rect 3608 440 3660 446
rect 3608 382 3660 388
rect 3690 417 3736 3511
rect 3769 3464 3815 3600
rect 3848 3545 3894 3557
rect 3848 3511 3854 3545
rect 3888 3511 3894 3545
rect 3690 383 3696 417
rect 3730 383 3736 417
rect 3690 100 3736 383
rect 3769 188 3815 464
rect 3769 151 3775 188
rect 3809 151 3815 188
rect 3769 139 3815 151
rect 3848 417 3894 3511
rect 4006 3545 4052 3557
rect 4006 3511 4012 3545
rect 4046 3511 4052 3545
rect 3927 446 3973 464
rect 3848 383 3854 417
rect 3888 383 3894 417
rect 3848 100 3894 383
rect 3924 440 3976 446
rect 3924 382 3976 388
rect 4006 417 4052 3511
rect 4085 3464 4131 3600
rect 4164 3545 4210 3557
rect 4164 3511 4170 3545
rect 4204 3511 4210 3545
rect 4006 383 4012 417
rect 4046 383 4052 417
rect 4006 100 4052 383
rect 4164 417 4210 3511
rect 4322 3545 4368 3557
rect 4322 3511 4328 3545
rect 4362 3511 4368 3545
rect 4243 446 4289 464
rect 4164 383 4170 417
rect 4204 383 4210 417
rect 4164 100 4210 383
rect 4240 440 4292 446
rect 4240 382 4292 388
rect 4322 417 4368 3511
rect 4401 3464 4447 3600
rect 4480 3545 4526 3557
rect 4480 3511 4486 3545
rect 4520 3511 4526 3545
rect 4322 383 4328 417
rect 4362 383 4368 417
rect 4322 100 4368 383
rect 4480 417 4526 3511
rect 4638 3545 4684 3557
rect 4638 3511 4644 3545
rect 4678 3511 4684 3545
rect 4559 446 4605 464
rect 4480 383 4486 417
rect 4520 383 4526 417
rect 4480 100 4526 383
rect 4556 440 4608 446
rect 4556 382 4608 388
rect 4638 417 4684 3511
rect 4717 3464 4763 3600
rect 4796 3545 4842 3557
rect 4796 3511 4802 3545
rect 4836 3511 4842 3545
rect 4638 383 4644 417
rect 4678 383 4684 417
rect 4638 100 4684 383
rect 4796 417 4842 3511
rect 4954 3545 5000 3557
rect 4954 3511 4960 3545
rect 4994 3511 5000 3545
rect 4875 446 4921 464
rect 4796 383 4802 417
rect 4836 383 4842 417
rect 4796 100 4842 383
rect 4872 440 4924 446
rect 4872 382 4924 388
rect 4954 417 5000 3511
rect 5033 3464 5079 3600
rect 5112 3545 5158 3557
rect 5112 3511 5118 3545
rect 5152 3511 5158 3545
rect 4954 383 4960 417
rect 4994 383 5000 417
rect 4954 100 5000 383
rect 5033 188 5079 464
rect 5033 151 5039 188
rect 5073 151 5079 188
rect 5033 139 5079 151
rect 5112 417 5158 3511
rect 5270 3545 5316 3557
rect 5270 3511 5276 3545
rect 5310 3511 5316 3545
rect 5191 446 5237 464
rect 5112 383 5118 417
rect 5152 383 5158 417
rect 5112 100 5158 383
rect 5188 440 5240 446
rect 5188 382 5240 388
rect 5270 417 5316 3511
rect 5349 3464 5395 3600
rect 5428 3545 5474 3557
rect 5428 3511 5434 3545
rect 5468 3511 5474 3545
rect 5270 383 5276 417
rect 5310 383 5316 417
rect 5270 100 5316 383
rect 5428 417 5474 3511
rect 5586 3545 5632 3557
rect 5586 3511 5592 3545
rect 5626 3511 5632 3545
rect 5507 446 5553 464
rect 5428 383 5434 417
rect 5468 383 5474 417
rect 5428 100 5474 383
rect 5504 440 5556 446
rect 5504 382 5556 388
rect 5586 417 5632 3511
rect 5665 3464 5711 3600
rect 5744 3545 5790 3557
rect 5744 3511 5750 3545
rect 5784 3511 5790 3545
rect 5586 383 5592 417
rect 5626 383 5632 417
rect 5586 100 5632 383
rect 5744 417 5790 3511
rect 5902 3545 5948 3557
rect 5902 3511 5908 3545
rect 5942 3511 5948 3545
rect 5823 446 5869 464
rect 5744 383 5750 417
rect 5784 383 5790 417
rect 5744 100 5790 383
rect 5820 440 5872 446
rect 5820 382 5872 388
rect 5902 417 5948 3511
rect 5981 3464 6027 3600
rect 6060 3545 6106 3557
rect 6060 3511 6066 3545
rect 6100 3511 6106 3545
rect 5902 383 5908 417
rect 5942 383 5948 417
rect 5902 100 5948 383
rect 6060 417 6106 3511
rect 6218 3545 6264 3557
rect 6218 3511 6224 3545
rect 6258 3511 6264 3545
rect 6139 446 6185 464
rect 6060 383 6066 417
rect 6100 383 6106 417
rect 6060 100 6106 383
rect 6136 440 6188 446
rect 6136 382 6188 388
rect 6218 417 6264 3511
rect 6297 3464 6343 3600
rect 6376 3545 6422 3557
rect 6376 3511 6382 3545
rect 6416 3511 6422 3545
rect 6218 383 6224 417
rect 6258 383 6264 417
rect 6218 100 6264 383
rect 6297 188 6343 464
rect 6297 151 6303 188
rect 6337 151 6343 188
rect 6297 139 6343 151
rect 6376 417 6422 3511
rect 6534 3545 6580 3557
rect 6534 3511 6540 3545
rect 6574 3511 6580 3545
rect 6455 446 6501 464
rect 6376 383 6382 417
rect 6416 383 6422 417
rect 6376 100 6422 383
rect 6452 440 6504 446
rect 6452 382 6504 388
rect 6534 417 6580 3511
rect 6613 3464 6659 3600
rect 6692 3545 6738 3557
rect 6692 3511 6698 3545
rect 6732 3511 6738 3545
rect 6534 383 6540 417
rect 6574 383 6580 417
rect 6534 100 6580 383
rect 6692 417 6738 3511
rect 6850 3545 6896 3557
rect 6850 3511 6856 3545
rect 6890 3511 6896 3545
rect 6771 446 6817 464
rect 6692 383 6698 417
rect 6732 383 6738 417
rect 6692 100 6738 383
rect 6768 440 6820 446
rect 6768 382 6820 388
rect 6850 417 6896 3511
rect 6929 3464 6975 3600
rect 6850 383 6856 417
rect 6890 383 6896 417
rect 6850 100 6896 383
rect 7400 124 7424 3600
rect 7476 3600 7600 3876
rect 7476 124 7500 3600
rect 7400 100 7500 124
rect -2472 80 6896 100
rect -2472 -80 -2426 80
rect 6060 -80 6896 80
rect -2472 -100 6896 -80
rect -2630 -417 -2624 -383
rect -2590 -417 -2584 -383
rect -2709 -455 -2663 -437
rect -2788 -1927 -2782 -1893
rect -2748 -1927 -2742 -1893
rect -2788 -1939 -2742 -1927
rect -2630 -1893 -2584 -417
rect -2551 -152 -2505 -140
rect -2551 -190 -2545 -152
rect -2511 -190 -2505 -152
rect -2551 -455 -2505 -190
rect -2472 -383 -2426 -100
rect -2472 -417 -2466 -383
rect -2432 -417 -2426 -383
rect -2630 -1927 -2624 -1893
rect -2590 -1927 -2584 -1893
rect -2630 -1939 -2584 -1927
rect -2551 -2000 -2505 -1855
rect -2472 -1893 -2426 -417
rect -2396 -379 -2344 -373
rect -2396 -437 -2344 -431
rect -2314 -383 -2268 -100
rect -2314 -417 -2308 -383
rect -2274 -417 -2268 -383
rect -2393 -455 -2347 -437
rect -2472 -1927 -2466 -1893
rect -2432 -1927 -2426 -1893
rect -2472 -1939 -2426 -1927
rect -2314 -1893 -2268 -417
rect -2156 -383 -2110 -100
rect -2156 -417 -2150 -383
rect -2116 -417 -2110 -383
rect -2314 -1927 -2308 -1893
rect -2274 -1927 -2268 -1893
rect -2314 -1939 -2268 -1927
rect -2235 -2000 -2189 -1855
rect -2156 -1893 -2110 -417
rect -2080 -379 -2028 -373
rect -2080 -437 -2028 -431
rect -1998 -383 -1952 -100
rect -1998 -417 -1992 -383
rect -1958 -417 -1952 -383
rect -2077 -455 -2031 -437
rect -2156 -1927 -2150 -1893
rect -2116 -1927 -2110 -1893
rect -2156 -1939 -2110 -1927
rect -1998 -1893 -1952 -417
rect -1840 -383 -1794 -100
rect -1840 -417 -1834 -383
rect -1800 -417 -1794 -383
rect -1998 -1927 -1992 -1893
rect -1958 -1927 -1952 -1893
rect -1998 -1939 -1952 -1927
rect -1919 -2000 -1873 -1855
rect -1840 -1893 -1794 -417
rect -1764 -379 -1712 -373
rect -1764 -437 -1712 -431
rect -1682 -383 -1636 -100
rect -1682 -417 -1676 -383
rect -1642 -417 -1636 -383
rect -1761 -455 -1715 -437
rect -1840 -1927 -1834 -1893
rect -1800 -1927 -1794 -1893
rect -1840 -1939 -1794 -1927
rect -1682 -1893 -1636 -417
rect -1524 -383 -1478 -100
rect -1524 -417 -1518 -383
rect -1484 -417 -1478 -383
rect -1682 -1927 -1676 -1893
rect -1642 -1927 -1636 -1893
rect -1682 -1939 -1636 -1927
rect -1603 -2000 -1557 -1855
rect -1524 -1893 -1478 -417
rect -1448 -379 -1396 -373
rect -1448 -437 -1396 -431
rect -1366 -383 -1320 -100
rect -1366 -417 -1360 -383
rect -1326 -417 -1320 -383
rect -1445 -455 -1399 -437
rect -1524 -1927 -1518 -1893
rect -1484 -1927 -1478 -1893
rect -1524 -1939 -1478 -1927
rect -1366 -1893 -1320 -417
rect -1287 -152 -1241 -140
rect -1287 -190 -1281 -152
rect -1247 -190 -1241 -152
rect -1287 -455 -1241 -190
rect -1208 -383 -1162 -100
rect -1208 -417 -1202 -383
rect -1168 -417 -1162 -383
rect -1366 -1927 -1360 -1893
rect -1326 -1927 -1320 -1893
rect -1366 -1939 -1320 -1927
rect -1287 -2000 -1241 -1855
rect -1208 -1893 -1162 -417
rect -1132 -379 -1080 -373
rect -1132 -437 -1080 -431
rect -1050 -383 -1004 -100
rect -1050 -417 -1044 -383
rect -1010 -417 -1004 -383
rect -1129 -455 -1083 -437
rect -1208 -1927 -1202 -1893
rect -1168 -1927 -1162 -1893
rect -1208 -1939 -1162 -1927
rect -1050 -1893 -1004 -417
rect -892 -383 -846 -100
rect -892 -417 -886 -383
rect -852 -417 -846 -383
rect -1050 -1927 -1044 -1893
rect -1010 -1927 -1004 -1893
rect -1050 -1939 -1004 -1927
rect -971 -2000 -925 -1855
rect -892 -1893 -846 -417
rect -816 -379 -764 -373
rect -816 -437 -764 -431
rect -734 -383 -688 -100
rect -734 -417 -728 -383
rect -694 -417 -688 -383
rect -813 -455 -767 -437
rect -892 -1927 -886 -1893
rect -852 -1927 -846 -1893
rect -892 -1939 -846 -1927
rect -734 -1893 -688 -417
rect -576 -383 -530 -100
rect -576 -417 -570 -383
rect -536 -417 -530 -383
rect -734 -1927 -728 -1893
rect -694 -1927 -688 -1893
rect -734 -1939 -688 -1927
rect -655 -2000 -609 -1855
rect -576 -1893 -530 -417
rect -500 -379 -448 -373
rect -500 -437 -448 -431
rect -418 -383 -372 -100
rect -418 -417 -412 -383
rect -378 -417 -372 -383
rect -497 -455 -451 -437
rect -576 -1927 -570 -1893
rect -536 -1927 -530 -1893
rect -576 -1939 -530 -1927
rect -418 -1893 -372 -417
rect -260 -383 -214 -100
rect -260 -417 -254 -383
rect -220 -417 -214 -383
rect -418 -1927 -412 -1893
rect -378 -1927 -372 -1893
rect -418 -1939 -372 -1927
rect -339 -2000 -293 -1855
rect -260 -1893 -214 -417
rect -184 -379 -132 -373
rect -184 -437 -132 -431
rect -102 -383 -56 -100
rect -102 -417 -96 -383
rect -62 -417 -56 -383
rect -181 -455 -135 -437
rect -260 -1927 -254 -1893
rect -220 -1927 -214 -1893
rect -260 -1939 -214 -1927
rect -102 -1893 -56 -417
rect -23 -152 23 -140
rect -23 -190 -17 -152
rect 17 -190 23 -152
rect -23 -455 23 -190
rect 56 -383 102 -100
rect 56 -417 62 -383
rect 96 -417 102 -383
rect -102 -1927 -96 -1893
rect -62 -1927 -56 -1893
rect -102 -1939 -56 -1927
rect -23 -2000 23 -1855
rect 56 -1893 102 -417
rect 132 -379 184 -373
rect 132 -437 184 -431
rect 214 -383 260 -100
rect 214 -417 220 -383
rect 254 -417 260 -383
rect 135 -455 181 -437
rect 56 -1927 62 -1893
rect 96 -1927 102 -1893
rect 56 -1939 102 -1927
rect 214 -1893 260 -417
rect 372 -383 418 -100
rect 372 -417 378 -383
rect 412 -417 418 -383
rect 214 -1927 220 -1893
rect 254 -1927 260 -1893
rect 214 -1939 260 -1927
rect 293 -2000 339 -1855
rect 372 -1893 418 -417
rect 448 -379 500 -373
rect 448 -437 500 -431
rect 530 -383 576 -100
rect 530 -417 536 -383
rect 570 -417 576 -383
rect 451 -455 497 -437
rect 372 -1927 378 -1893
rect 412 -1927 418 -1893
rect 372 -1939 418 -1927
rect 530 -1893 576 -417
rect 688 -383 734 -100
rect 688 -417 694 -383
rect 728 -417 734 -383
rect 530 -1927 536 -1893
rect 570 -1927 576 -1893
rect 530 -1939 576 -1927
rect 609 -2000 655 -1855
rect 688 -1893 734 -417
rect 764 -379 816 -373
rect 764 -437 816 -431
rect 846 -383 892 -100
rect 846 -417 852 -383
rect 886 -417 892 -383
rect 767 -455 813 -437
rect 688 -1927 694 -1893
rect 728 -1927 734 -1893
rect 688 -1939 734 -1927
rect 846 -1893 892 -417
rect 1004 -383 1050 -100
rect 1004 -417 1010 -383
rect 1044 -417 1050 -383
rect 846 -1927 852 -1893
rect 886 -1927 892 -1893
rect 846 -1939 892 -1927
rect 925 -2000 971 -1855
rect 1004 -1893 1050 -417
rect 1080 -379 1132 -373
rect 1080 -437 1132 -431
rect 1162 -383 1208 -100
rect 1162 -417 1168 -383
rect 1202 -417 1208 -383
rect 1083 -455 1129 -437
rect 1004 -1927 1010 -1893
rect 1044 -1927 1050 -1893
rect 1004 -1939 1050 -1927
rect 1162 -1893 1208 -417
rect 1241 -152 1287 -140
rect 1241 -190 1247 -152
rect 1281 -190 1287 -152
rect 1241 -455 1287 -190
rect 1320 -383 1366 -100
rect 1320 -417 1326 -383
rect 1360 -417 1366 -383
rect 1162 -1927 1168 -1893
rect 1202 -1927 1208 -1893
rect 1162 -1939 1208 -1927
rect 1241 -2000 1287 -1855
rect 1320 -1893 1366 -417
rect 1396 -379 1448 -373
rect 1396 -437 1448 -431
rect 1478 -383 1524 -100
rect 1478 -417 1484 -383
rect 1518 -417 1524 -383
rect 1399 -455 1445 -437
rect 1320 -1927 1326 -1893
rect 1360 -1927 1366 -1893
rect 1320 -1939 1366 -1927
rect 1478 -1893 1524 -417
rect 1636 -383 1682 -100
rect 1636 -417 1642 -383
rect 1676 -417 1682 -383
rect 1478 -1927 1484 -1893
rect 1518 -1927 1524 -1893
rect 1478 -1939 1524 -1927
rect 1557 -2000 1603 -1855
rect 1636 -1893 1682 -417
rect 1712 -379 1764 -373
rect 1712 -437 1764 -431
rect 1794 -383 1840 -100
rect 1794 -417 1800 -383
rect 1834 -417 1840 -383
rect 1715 -455 1761 -437
rect 1636 -1927 1642 -1893
rect 1676 -1927 1682 -1893
rect 1636 -1939 1682 -1927
rect 1794 -1893 1840 -417
rect 1952 -383 1998 -100
rect 1952 -417 1958 -383
rect 1992 -417 1998 -383
rect 1794 -1927 1800 -1893
rect 1834 -1927 1840 -1893
rect 1794 -1939 1840 -1927
rect 1873 -2000 1919 -1855
rect 1952 -1893 1998 -417
rect 2028 -379 2080 -373
rect 2028 -437 2080 -431
rect 2110 -383 2156 -100
rect 2110 -417 2116 -383
rect 2150 -417 2156 -383
rect 2031 -455 2077 -437
rect 1952 -1927 1958 -1893
rect 1992 -1927 1998 -1893
rect 1952 -1939 1998 -1927
rect 2110 -1893 2156 -417
rect 2268 -383 2314 -100
rect 2268 -417 2274 -383
rect 2308 -417 2314 -383
rect 2110 -1927 2116 -1893
rect 2150 -1927 2156 -1893
rect 2110 -1939 2156 -1927
rect 2189 -2000 2235 -1855
rect 2268 -1893 2314 -417
rect 2344 -379 2396 -373
rect 2344 -437 2396 -431
rect 2426 -383 2472 -100
rect 2426 -417 2432 -383
rect 2466 -417 2472 -383
rect 2347 -455 2393 -437
rect 2268 -1927 2274 -1893
rect 2308 -1927 2314 -1893
rect 2268 -1939 2314 -1927
rect 2426 -1893 2472 -417
rect 2505 -152 2551 -140
rect 2505 -190 2511 -152
rect 2545 -190 2551 -152
rect 2505 -455 2551 -190
rect 2584 -383 2630 -100
rect 2584 -417 2590 -383
rect 2624 -417 2630 -383
rect 2426 -1927 2432 -1893
rect 2466 -1927 2472 -1893
rect 2426 -1939 2472 -1927
rect 2505 -2000 2551 -1855
rect 2584 -1893 2630 -417
rect 2660 -379 2712 -373
rect 2660 -437 2712 -431
rect 2742 -383 2788 -100
rect 2742 -417 2748 -383
rect 2782 -417 2788 -383
rect 2663 -455 2709 -437
rect 2584 -1927 2590 -1893
rect 2624 -1927 2630 -1893
rect 2584 -1939 2630 -1927
rect 2742 -1893 2788 -417
rect 2900 -383 2946 -100
rect 2900 -417 2906 -383
rect 2940 -417 2946 -383
rect 2742 -1927 2748 -1893
rect 2782 -1927 2788 -1893
rect 2742 -1939 2788 -1927
rect 2821 -2000 2867 -1855
rect 2900 -1893 2946 -417
rect 2976 -379 3028 -373
rect 2976 -437 3028 -431
rect 3058 -383 3104 -100
rect 3058 -417 3064 -383
rect 3098 -417 3104 -383
rect 2979 -455 3025 -437
rect 2900 -1927 2906 -1893
rect 2940 -1927 2946 -1893
rect 2900 -1939 2946 -1927
rect 3058 -1893 3104 -417
rect 3216 -383 3262 -100
rect 3216 -417 3222 -383
rect 3256 -417 3262 -383
rect 3058 -1927 3064 -1893
rect 3098 -1927 3104 -1893
rect 3058 -1939 3104 -1927
rect 3137 -2000 3183 -1855
rect 3216 -1893 3262 -417
rect 3292 -379 3344 -373
rect 3292 -437 3344 -431
rect 3374 -383 3420 -100
rect 3374 -417 3380 -383
rect 3414 -417 3420 -383
rect 3295 -455 3341 -437
rect 3216 -1927 3222 -1893
rect 3256 -1927 3262 -1893
rect 3216 -1939 3262 -1927
rect 3374 -1893 3420 -417
rect 3532 -383 3578 -100
rect 3532 -417 3538 -383
rect 3572 -417 3578 -383
rect 3374 -1927 3380 -1893
rect 3414 -1927 3420 -1893
rect 3374 -1939 3420 -1927
rect 3453 -2000 3499 -1855
rect 3532 -1893 3578 -417
rect 3608 -379 3660 -373
rect 3608 -437 3660 -431
rect 3690 -383 3736 -100
rect 3690 -417 3696 -383
rect 3730 -417 3736 -383
rect 3611 -455 3657 -437
rect 3532 -1927 3538 -1893
rect 3572 -1927 3578 -1893
rect 3532 -1939 3578 -1927
rect 3690 -1893 3736 -417
rect 3769 -152 3815 -140
rect 3769 -190 3775 -152
rect 3809 -190 3815 -152
rect 3769 -455 3815 -190
rect 3848 -383 3894 -100
rect 3848 -417 3854 -383
rect 3888 -417 3894 -383
rect 3690 -1927 3696 -1893
rect 3730 -1927 3736 -1893
rect 3690 -1939 3736 -1927
rect 3769 -2000 3815 -1855
rect 3848 -1893 3894 -417
rect 3924 -379 3976 -373
rect 3924 -437 3976 -431
rect 4006 -383 4052 -100
rect 4006 -417 4012 -383
rect 4046 -417 4052 -383
rect 3927 -455 3973 -437
rect 3848 -1927 3854 -1893
rect 3888 -1927 3894 -1893
rect 3848 -1939 3894 -1927
rect 4006 -1893 4052 -417
rect 4164 -383 4210 -100
rect 4164 -417 4170 -383
rect 4204 -417 4210 -383
rect 4006 -1927 4012 -1893
rect 4046 -1927 4052 -1893
rect 4006 -1939 4052 -1927
rect 4085 -2000 4131 -1855
rect 4164 -1893 4210 -417
rect 4240 -379 4292 -373
rect 4240 -437 4292 -431
rect 4322 -383 4368 -100
rect 4322 -417 4328 -383
rect 4362 -417 4368 -383
rect 4243 -455 4289 -437
rect 4164 -1927 4170 -1893
rect 4204 -1927 4210 -1893
rect 4164 -1939 4210 -1927
rect 4322 -1893 4368 -417
rect 4480 -383 4526 -100
rect 4480 -417 4486 -383
rect 4520 -417 4526 -383
rect 4322 -1927 4328 -1893
rect 4362 -1927 4368 -1893
rect 4322 -1939 4368 -1927
rect 4401 -2000 4447 -1855
rect 4480 -1893 4526 -417
rect 4556 -379 4608 -373
rect 4556 -437 4608 -431
rect 4638 -383 4684 -100
rect 4638 -417 4644 -383
rect 4678 -417 4684 -383
rect 4559 -455 4605 -437
rect 4480 -1927 4486 -1893
rect 4520 -1927 4526 -1893
rect 4480 -1939 4526 -1927
rect 4638 -1893 4684 -417
rect 4796 -383 4842 -100
rect 4796 -417 4802 -383
rect 4836 -417 4842 -383
rect 4638 -1927 4644 -1893
rect 4678 -1927 4684 -1893
rect 4638 -1939 4684 -1927
rect 4717 -2000 4763 -1855
rect 4796 -1893 4842 -417
rect 4872 -379 4924 -373
rect 4872 -437 4924 -431
rect 4954 -383 5000 -100
rect 4954 -417 4960 -383
rect 4994 -417 5000 -383
rect 4875 -455 4921 -437
rect 4796 -1927 4802 -1893
rect 4836 -1927 4842 -1893
rect 4796 -1939 4842 -1927
rect 4954 -1893 5000 -417
rect 5033 -152 5079 -140
rect 5033 -190 5039 -152
rect 5073 -190 5079 -152
rect 5033 -455 5079 -190
rect 5112 -383 5158 -100
rect 5112 -417 5118 -383
rect 5152 -417 5158 -383
rect 4954 -1927 4960 -1893
rect 4994 -1927 5000 -1893
rect 4954 -1939 5000 -1927
rect 5033 -2000 5079 -1855
rect 5112 -1893 5158 -417
rect 5188 -379 5240 -373
rect 5188 -437 5240 -431
rect 5270 -383 5316 -100
rect 5270 -417 5276 -383
rect 5310 -417 5316 -383
rect 5191 -455 5237 -437
rect 5112 -1927 5118 -1893
rect 5152 -1927 5158 -1893
rect 5112 -1939 5158 -1927
rect 5270 -1893 5316 -417
rect 5428 -383 5474 -100
rect 5428 -417 5434 -383
rect 5468 -417 5474 -383
rect 5270 -1927 5276 -1893
rect 5310 -1927 5316 -1893
rect 5270 -1939 5316 -1927
rect 5349 -2000 5395 -1855
rect 5428 -1893 5474 -417
rect 5504 -379 5556 -373
rect 5504 -437 5556 -431
rect 5586 -383 5632 -100
rect 5586 -417 5592 -383
rect 5626 -417 5632 -383
rect 5507 -455 5553 -437
rect 5428 -1927 5434 -1893
rect 5468 -1927 5474 -1893
rect 5428 -1939 5474 -1927
rect 5586 -1893 5632 -417
rect 5744 -383 5790 -100
rect 5744 -417 5750 -383
rect 5784 -417 5790 -383
rect 5586 -1927 5592 -1893
rect 5626 -1927 5632 -1893
rect 5586 -1939 5632 -1927
rect 5665 -2000 5711 -1855
rect 5744 -1893 5790 -417
rect 5820 -379 5872 -373
rect 5820 -437 5872 -431
rect 5902 -383 5948 -100
rect 5902 -417 5908 -383
rect 5942 -417 5948 -383
rect 5823 -455 5869 -437
rect 5744 -1927 5750 -1893
rect 5784 -1927 5790 -1893
rect 5744 -1939 5790 -1927
rect 5902 -1893 5948 -417
rect 6060 -383 6106 -100
rect 6060 -417 6066 -383
rect 6100 -417 6106 -383
rect 5902 -1927 5908 -1893
rect 5942 -1927 5948 -1893
rect 5902 -1939 5948 -1927
rect 5981 -2000 6027 -1855
rect 6060 -1893 6106 -417
rect 6136 -379 6188 -373
rect 6136 -437 6188 -431
rect 6218 -383 6264 -100
rect 6218 -417 6224 -383
rect 6258 -417 6264 -383
rect 6139 -455 6185 -437
rect 6060 -1927 6066 -1893
rect 6100 -1927 6106 -1893
rect 6060 -1939 6106 -1927
rect 6218 -1893 6264 -417
rect 6297 -152 6343 -140
rect 6297 -190 6303 -152
rect 6337 -190 6343 -152
rect 6297 -455 6343 -190
rect 6376 -383 6422 -100
rect 6376 -417 6382 -383
rect 6416 -417 6422 -383
rect 6218 -1927 6224 -1893
rect 6258 -1927 6264 -1893
rect 6218 -1939 6264 -1927
rect 6297 -2000 6343 -1855
rect 6376 -1893 6422 -417
rect 6452 -379 6504 -373
rect 6452 -437 6504 -431
rect 6534 -383 6580 -100
rect 6534 -417 6540 -383
rect 6574 -417 6580 -383
rect 6455 -455 6501 -437
rect 6376 -1927 6382 -1893
rect 6416 -1927 6422 -1893
rect 6376 -1939 6422 -1927
rect 6534 -1893 6580 -417
rect 6692 -383 6738 -100
rect 6692 -417 6698 -383
rect 6732 -417 6738 -383
rect 6534 -1927 6540 -1893
rect 6574 -1927 6580 -1893
rect 6534 -1939 6580 -1927
rect 6613 -2000 6659 -1855
rect 6692 -1893 6738 -417
rect 6768 -379 6820 -373
rect 6768 -437 6820 -431
rect 6850 -383 6896 -100
rect 6850 -417 6856 -383
rect 6890 -417 6896 -383
rect 6771 -455 6817 -437
rect 6692 -1927 6698 -1893
rect 6732 -1927 6738 -1893
rect 6692 -1939 6738 -1927
rect 6850 -1893 6896 -417
rect 7400 -124 7500 -100
rect 6850 -1927 6856 -1893
rect 6890 -1927 6896 -1893
rect 6850 -1939 6896 -1927
rect 6929 -2000 6975 -1855
rect 7400 -2000 7424 -124
rect -8324 -2224 7424 -2000
rect 7476 -2000 7500 -124
rect 7476 -2276 7600 -2000
rect -8500 -2400 7600 -2276
<< via1 >>
rect -6820 388 -6768 440
rect -7739 -943 -7682 -907
rect -7739 -959 -7682 -943
rect -7423 -943 -7366 -907
rect -7423 -959 -7366 -943
rect -6820 -431 -6768 -379
rect -6504 388 -6452 440
rect -6188 388 -6136 440
rect -5872 388 -5820 440
rect -6560 -80 -6246 80
rect -6504 -431 -6452 -379
rect -6188 -431 -6136 -379
rect -5872 -431 -5820 -379
rect -5556 388 -5504 440
rect -5240 388 -5188 440
rect -4924 388 -4872 440
rect -4608 388 -4556 440
rect -4292 388 -4240 440
rect -3976 388 -3924 440
rect -3660 388 -3608 440
rect -3344 388 -3292 440
rect -3028 388 -2976 440
rect -2712 388 -2660 440
rect -5562 -80 -3078 80
rect -5556 -431 -5504 -379
rect -5240 -431 -5188 -379
rect -4924 -431 -4872 -379
rect -4608 -431 -4556 -379
rect -4292 -431 -4240 -379
rect -3976 -431 -3924 -379
rect -3660 -431 -3608 -379
rect -3344 -431 -3292 -379
rect -3028 -431 -2976 -379
rect -2712 -431 -2660 -379
rect -2396 388 -2344 440
rect -2080 388 -2028 440
rect -1764 388 -1712 440
rect -1448 388 -1396 440
rect -1132 388 -1080 440
rect -816 388 -764 440
rect -500 388 -448 440
rect -184 388 -132 440
rect 132 388 184 440
rect 448 388 500 440
rect 764 388 816 440
rect 1080 388 1132 440
rect 1396 388 1448 440
rect 1712 388 1764 440
rect 2028 388 2080 440
rect 2344 388 2396 440
rect 2660 388 2712 440
rect 2976 388 3028 440
rect 3292 388 3344 440
rect 3608 388 3660 440
rect 3924 388 3976 440
rect 4240 388 4292 440
rect 4556 388 4608 440
rect 4872 388 4924 440
rect 5188 388 5240 440
rect 5504 388 5556 440
rect 5820 388 5872 440
rect 6136 388 6188 440
rect 6452 388 6504 440
rect 6768 388 6820 440
rect -2426 -80 6060 80
rect -2396 -431 -2344 -379
rect -2080 -431 -2028 -379
rect -1764 -431 -1712 -379
rect -1448 -431 -1396 -379
rect -1132 -431 -1080 -379
rect -816 -431 -764 -379
rect -500 -431 -448 -379
rect -184 -431 -132 -379
rect 132 -431 184 -379
rect 448 -431 500 -379
rect 764 -431 816 -379
rect 1080 -431 1132 -379
rect 1396 -431 1448 -379
rect 1712 -431 1764 -379
rect 2028 -431 2080 -379
rect 2344 -431 2396 -379
rect 2660 -431 2712 -379
rect 2976 -431 3028 -379
rect 3292 -431 3344 -379
rect 3608 -431 3660 -379
rect 3924 -431 3976 -379
rect 4240 -431 4292 -379
rect 4556 -431 4608 -379
rect 4872 -431 4924 -379
rect 5188 -431 5240 -379
rect 5504 -431 5556 -379
rect 5820 -431 5872 -379
rect 6136 -431 6188 -379
rect 6452 -431 6504 -379
rect 6768 -431 6820 -379
<< metal2 >>
rect -6826 388 -6820 440
rect -6768 388 -6762 440
rect -6510 388 -6504 440
rect -6452 388 -6188 440
rect -6136 388 -5872 440
rect -5820 388 -5814 440
rect -6817 214 -6771 388
rect -6817 100 -6580 214
rect -6510 140 -5814 388
rect -5562 388 -5556 440
rect -5504 388 -5240 440
rect -5188 388 -4924 440
rect -4872 388 -4608 440
rect -4556 388 -4292 440
rect -4240 388 -3976 440
rect -3924 388 -3660 440
rect -3608 388 -3344 440
rect -3292 388 -3028 440
rect -2976 388 -2712 440
rect -2660 388 -2654 440
rect -5562 140 -2654 388
rect -2402 388 -2396 440
rect -2344 388 -2080 440
rect -2028 388 -1764 440
rect -1712 388 -1448 440
rect -1396 388 -1132 440
rect -1080 388 -816 440
rect -764 388 -500 440
rect -448 388 -184 440
rect -132 388 132 440
rect 184 388 448 440
rect 500 388 764 440
rect 816 388 1080 440
rect 1132 388 1396 440
rect 1448 388 1712 440
rect 1764 388 2028 440
rect 2080 388 2344 440
rect 2396 388 2660 440
rect 2712 388 2976 440
rect 3028 388 3292 440
rect 3344 388 3608 440
rect 3660 388 3924 440
rect 3976 388 4240 440
rect 4292 388 4556 440
rect 4608 388 4872 440
rect 4924 388 5188 440
rect 5240 388 5504 440
rect 5556 388 5820 440
rect 5872 388 6136 440
rect 6188 388 6452 440
rect 6504 388 6768 440
rect 6820 388 7500 440
rect -2402 140 7500 388
rect -6060 100 -5814 140
rect -2900 100 -2654 140
rect -6817 91 -6218 100
rect -6652 80 -6218 91
rect -6652 -80 -6560 80
rect -6246 -80 -6218 80
rect -6652 -91 -6218 -80
rect -6817 -100 -6218 -91
rect -6060 80 -3058 100
rect -6060 -80 -5562 80
rect -3078 -80 -3058 80
rect -6060 -100 -3058 -80
rect -2900 80 6106 100
rect -2900 -80 -2426 80
rect 6060 -80 6106 80
rect -2900 -100 6106 -80
rect -6817 -205 -6580 -100
rect -6060 -140 -5814 -100
rect -2900 -140 -2654 -100
rect 6163 -140 7500 140
rect -6817 -379 -6771 -205
rect -6510 -379 -5814 -140
rect -6826 -431 -6820 -379
rect -6768 -431 -6762 -379
rect -6510 -431 -6504 -379
rect -6452 -431 -6188 -379
rect -6136 -431 -5872 -379
rect -5820 -431 -5814 -379
rect -5562 -379 -2654 -140
rect -5562 -431 -5556 -379
rect -5504 -431 -5240 -379
rect -5188 -431 -4924 -379
rect -4872 -431 -4608 -379
rect -4556 -431 -4292 -379
rect -4240 -431 -3976 -379
rect -3924 -431 -3660 -379
rect -3608 -431 -3344 -379
rect -3292 -431 -3028 -379
rect -2976 -431 -2712 -379
rect -2660 -431 -2654 -379
rect -2402 -379 7500 -140
rect -2402 -431 -2396 -379
rect -2344 -431 -2080 -379
rect -2028 -431 -1764 -379
rect -1712 -431 -1448 -379
rect -1396 -431 -1132 -379
rect -1080 -431 -816 -379
rect -764 -431 -500 -379
rect -448 -431 -184 -379
rect -132 -431 132 -379
rect 184 -431 448 -379
rect 500 -431 764 -379
rect 816 -431 1080 -379
rect 1132 -431 1396 -379
rect 1448 -431 1712 -379
rect 1764 -431 2028 -379
rect 2080 -431 2344 -379
rect 2396 -431 2660 -379
rect 2712 -431 2976 -379
rect 3028 -431 3292 -379
rect 3344 -431 3608 -379
rect 3660 -431 3924 -379
rect 3976 -431 4240 -379
rect 4292 -431 4556 -379
rect 4608 -431 4872 -379
rect 4924 -431 5188 -379
rect 5240 -431 5504 -379
rect 5556 -431 5820 -379
rect 5872 -431 6136 -379
rect 6188 -431 6452 -379
rect 6504 -431 6768 -379
rect 6820 -431 7500 -379
rect -7739 -907 -7682 -897
rect -8012 -959 -7739 -934
rect -7423 -907 -7366 -897
rect -8012 -994 -7682 -959
rect -7483 -959 -7423 -934
rect -7483 -994 -7366 -959
rect -7483 -1038 -7423 -994
rect -8012 -1098 -7423 -1038
use sky130_fd_pr__pfet_g5v0d10v5_RTDP6L  xm4
timestamp 1624430562
transform 1 0 -7552 0 1 864
box -411 -500 411 500
use sky130_fd_pr__nfet_g5v0d10v5_3BH9ZH  xm3
timestamp 1624430562
transform 1 0 -7552 0 1 -655
box -345 -288 345 288
use sky130_fd_pr__pfet_g5v0d10v5_7WGKBW  xm2
timestamp 1624430562
transform 1 0 0 0 1 1964
box -7047 -1600 7047 1600
use sky130_fd_pr__nfet_g5v0d10v5_WQT6C6  xm1
timestamp 1624430562
transform 1 0 0 0 1 -1155
box -6981 -788 6981 788
<< labels >>
flabel metal2 7500 -431 7500 440 1 FreeSans 240 0 0 0 out
port 3 n
flabel metal1 -8500 3600 -8500 4000 3 FreeSans 240 0 0 0 vdd
port 4 e
flabel metal1 -8500 -2400 -8500 -2000 3 FreeSans 240 0 0 0 vss
port 5 e
flabel metal2 -8012 -994 -8012 -934 1 FreeSans 240 0 0 0 in_p
port 2 n
flabel metal2 -8012 -1098 -8012 -1038 1 FreeSans 240 0 0 0 in_m
port 1 n
<< end >>
