magic
tech sky130A
magscale 1 2
timestamp 1624430562
<< error_p >>
rect -6995 -500 -6937 500
rect -6737 -500 -6679 500
rect -6479 -500 -6421 500
rect -6221 -500 -6163 500
rect -5963 -500 -5905 500
rect -5705 -500 -5647 500
rect -5447 -500 -5389 500
rect -5189 -500 -5131 500
rect -4931 -500 -4873 500
rect -4673 -500 -4615 500
rect -4415 -500 -4357 500
rect -4157 -500 -4099 500
rect -3899 -500 -3841 500
rect -3641 -500 -3583 500
rect -3383 -500 -3325 500
rect -3125 -500 -3067 500
rect -2867 -500 -2809 500
rect -2609 -500 -2551 500
rect -2351 -500 -2293 500
rect -2093 -500 -2035 500
rect -1835 -500 -1777 500
rect -1577 -500 -1519 500
rect -1319 -500 -1261 500
rect -1061 -500 -1003 500
rect -803 -500 -745 500
rect -545 -500 -487 500
rect -287 -500 -229 500
rect -29 -500 29 500
rect 229 -500 287 500
rect 487 -500 545 500
rect 745 -500 803 500
rect 1003 -500 1061 500
rect 1261 -500 1319 500
rect 1519 -500 1577 500
rect 1777 -500 1835 500
rect 2035 -500 2093 500
rect 2293 -500 2351 500
rect 2551 -500 2609 500
rect 2809 -500 2867 500
rect 3067 -500 3125 500
rect 3325 -500 3383 500
rect 3583 -500 3641 500
rect 3841 -500 3899 500
rect 4099 -500 4157 500
rect 4357 -500 4415 500
rect 4615 -500 4673 500
rect 4873 -500 4931 500
rect 5131 -500 5189 500
rect 5389 -500 5447 500
rect 5647 -500 5705 500
rect 5905 -500 5963 500
rect 6163 -500 6221 500
rect 6421 -500 6479 500
rect 6679 -500 6737 500
rect 6937 -500 6995 500
<< mvnmos >>
rect -6937 -500 -6737 500
rect -6679 -500 -6479 500
rect -6421 -500 -6221 500
rect -6163 -500 -5963 500
rect -5905 -500 -5705 500
rect -5647 -500 -5447 500
rect -5389 -500 -5189 500
rect -5131 -500 -4931 500
rect -4873 -500 -4673 500
rect -4615 -500 -4415 500
rect -4357 -500 -4157 500
rect -4099 -500 -3899 500
rect -3841 -500 -3641 500
rect -3583 -500 -3383 500
rect -3325 -500 -3125 500
rect -3067 -500 -2867 500
rect -2809 -500 -2609 500
rect -2551 -500 -2351 500
rect -2293 -500 -2093 500
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
rect 2093 -500 2293 500
rect 2351 -500 2551 500
rect 2609 -500 2809 500
rect 2867 -500 3067 500
rect 3125 -500 3325 500
rect 3383 -500 3583 500
rect 3641 -500 3841 500
rect 3899 -500 4099 500
rect 4157 -500 4357 500
rect 4415 -500 4615 500
rect 4673 -500 4873 500
rect 4931 -500 5131 500
rect 5189 -500 5389 500
rect 5447 -500 5647 500
rect 5705 -500 5905 500
rect 5963 -500 6163 500
rect 6221 -500 6421 500
rect 6479 -500 6679 500
rect 6737 -500 6937 500
<< mvndiff >>
rect -6995 488 -6937 500
rect -6995 -488 -6983 488
rect -6949 -488 -6937 488
rect -6995 -500 -6937 -488
rect -6737 488 -6679 500
rect -6737 -488 -6725 488
rect -6691 -488 -6679 488
rect -6737 -500 -6679 -488
rect -6479 488 -6421 500
rect -6479 -488 -6467 488
rect -6433 -488 -6421 488
rect -6479 -500 -6421 -488
rect -6221 488 -6163 500
rect -6221 -488 -6209 488
rect -6175 -488 -6163 488
rect -6221 -500 -6163 -488
rect -5963 488 -5905 500
rect -5963 -488 -5951 488
rect -5917 -488 -5905 488
rect -5963 -500 -5905 -488
rect -5705 488 -5647 500
rect -5705 -488 -5693 488
rect -5659 -488 -5647 488
rect -5705 -500 -5647 -488
rect -5447 488 -5389 500
rect -5447 -488 -5435 488
rect -5401 -488 -5389 488
rect -5447 -500 -5389 -488
rect -5189 488 -5131 500
rect -5189 -488 -5177 488
rect -5143 -488 -5131 488
rect -5189 -500 -5131 -488
rect -4931 488 -4873 500
rect -4931 -488 -4919 488
rect -4885 -488 -4873 488
rect -4931 -500 -4873 -488
rect -4673 488 -4615 500
rect -4673 -488 -4661 488
rect -4627 -488 -4615 488
rect -4673 -500 -4615 -488
rect -4415 488 -4357 500
rect -4415 -488 -4403 488
rect -4369 -488 -4357 488
rect -4415 -500 -4357 -488
rect -4157 488 -4099 500
rect -4157 -488 -4145 488
rect -4111 -488 -4099 488
rect -4157 -500 -4099 -488
rect -3899 488 -3841 500
rect -3899 -488 -3887 488
rect -3853 -488 -3841 488
rect -3899 -500 -3841 -488
rect -3641 488 -3583 500
rect -3641 -488 -3629 488
rect -3595 -488 -3583 488
rect -3641 -500 -3583 -488
rect -3383 488 -3325 500
rect -3383 -488 -3371 488
rect -3337 -488 -3325 488
rect -3383 -500 -3325 -488
rect -3125 488 -3067 500
rect -3125 -488 -3113 488
rect -3079 -488 -3067 488
rect -3125 -500 -3067 -488
rect -2867 488 -2809 500
rect -2867 -488 -2855 488
rect -2821 -488 -2809 488
rect -2867 -500 -2809 -488
rect -2609 488 -2551 500
rect -2609 -488 -2597 488
rect -2563 -488 -2551 488
rect -2609 -500 -2551 -488
rect -2351 488 -2293 500
rect -2351 -488 -2339 488
rect -2305 -488 -2293 488
rect -2351 -500 -2293 -488
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
rect 2293 488 2351 500
rect 2293 -488 2305 488
rect 2339 -488 2351 488
rect 2293 -500 2351 -488
rect 2551 488 2609 500
rect 2551 -488 2563 488
rect 2597 -488 2609 488
rect 2551 -500 2609 -488
rect 2809 488 2867 500
rect 2809 -488 2821 488
rect 2855 -488 2867 488
rect 2809 -500 2867 -488
rect 3067 488 3125 500
rect 3067 -488 3079 488
rect 3113 -488 3125 488
rect 3067 -500 3125 -488
rect 3325 488 3383 500
rect 3325 -488 3337 488
rect 3371 -488 3383 488
rect 3325 -500 3383 -488
rect 3583 488 3641 500
rect 3583 -488 3595 488
rect 3629 -488 3641 488
rect 3583 -500 3641 -488
rect 3841 488 3899 500
rect 3841 -488 3853 488
rect 3887 -488 3899 488
rect 3841 -500 3899 -488
rect 4099 488 4157 500
rect 4099 -488 4111 488
rect 4145 -488 4157 488
rect 4099 -500 4157 -488
rect 4357 488 4415 500
rect 4357 -488 4369 488
rect 4403 -488 4415 488
rect 4357 -500 4415 -488
rect 4615 488 4673 500
rect 4615 -488 4627 488
rect 4661 -488 4673 488
rect 4615 -500 4673 -488
rect 4873 488 4931 500
rect 4873 -488 4885 488
rect 4919 -488 4931 488
rect 4873 -500 4931 -488
rect 5131 488 5189 500
rect 5131 -488 5143 488
rect 5177 -488 5189 488
rect 5131 -500 5189 -488
rect 5389 488 5447 500
rect 5389 -488 5401 488
rect 5435 -488 5447 488
rect 5389 -500 5447 -488
rect 5647 488 5705 500
rect 5647 -488 5659 488
rect 5693 -488 5705 488
rect 5647 -500 5705 -488
rect 5905 488 5963 500
rect 5905 -488 5917 488
rect 5951 -488 5963 488
rect 5905 -500 5963 -488
rect 6163 488 6221 500
rect 6163 -488 6175 488
rect 6209 -488 6221 488
rect 6163 -500 6221 -488
rect 6421 488 6479 500
rect 6421 -488 6433 488
rect 6467 -488 6479 488
rect 6421 -500 6479 -488
rect 6679 488 6737 500
rect 6679 -488 6691 488
rect 6725 -488 6737 488
rect 6679 -500 6737 -488
rect 6937 488 6995 500
rect 6937 -488 6949 488
rect 6983 -488 6995 488
rect 6937 -500 6995 -488
<< mvndiffc >>
rect -6983 -488 -6949 488
rect -6725 -488 -6691 488
rect -6467 -488 -6433 488
rect -6209 -488 -6175 488
rect -5951 -488 -5917 488
rect -5693 -488 -5659 488
rect -5435 -488 -5401 488
rect -5177 -488 -5143 488
rect -4919 -488 -4885 488
rect -4661 -488 -4627 488
rect -4403 -488 -4369 488
rect -4145 -488 -4111 488
rect -3887 -488 -3853 488
rect -3629 -488 -3595 488
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect 3595 -488 3629 488
rect 3853 -488 3887 488
rect 4111 -488 4145 488
rect 4369 -488 4403 488
rect 4627 -488 4661 488
rect 4885 -488 4919 488
rect 5143 -488 5177 488
rect 5401 -488 5435 488
rect 5659 -488 5693 488
rect 5917 -488 5951 488
rect 6175 -488 6209 488
rect 6433 -488 6467 488
rect 6691 -488 6725 488
rect 6949 -488 6983 488
<< poly >>
rect -6903 572 -6771 588
rect -6903 555 -6887 572
rect -6937 538 -6887 555
rect -6787 555 -6771 572
rect -6645 572 -6513 588
rect -6645 555 -6629 572
rect -6787 538 -6737 555
rect -6937 500 -6737 538
rect -6679 538 -6629 555
rect -6529 555 -6513 572
rect -6387 572 -6255 588
rect -6387 555 -6371 572
rect -6529 538 -6479 555
rect -6679 500 -6479 538
rect -6421 538 -6371 555
rect -6271 555 -6255 572
rect -6129 572 -5997 588
rect -6129 555 -6113 572
rect -6271 538 -6221 555
rect -6421 500 -6221 538
rect -6163 538 -6113 555
rect -6013 555 -5997 572
rect -5871 572 -5739 588
rect -5871 555 -5855 572
rect -6013 538 -5963 555
rect -6163 500 -5963 538
rect -5905 538 -5855 555
rect -5755 555 -5739 572
rect -5613 572 -5481 588
rect -5613 555 -5597 572
rect -5755 538 -5705 555
rect -5905 500 -5705 538
rect -5647 538 -5597 555
rect -5497 555 -5481 572
rect -5355 572 -5223 588
rect -5355 555 -5339 572
rect -5497 538 -5447 555
rect -5647 500 -5447 538
rect -5389 538 -5339 555
rect -5239 555 -5223 572
rect -5097 572 -4965 588
rect -5097 555 -5081 572
rect -5239 538 -5189 555
rect -5389 500 -5189 538
rect -5131 538 -5081 555
rect -4981 555 -4965 572
rect -4839 572 -4707 588
rect -4839 555 -4823 572
rect -4981 538 -4931 555
rect -5131 500 -4931 538
rect -4873 538 -4823 555
rect -4723 555 -4707 572
rect -4581 572 -4449 588
rect -4581 555 -4565 572
rect -4723 538 -4673 555
rect -4873 500 -4673 538
rect -4615 538 -4565 555
rect -4465 555 -4449 572
rect -4323 572 -4191 588
rect -4323 555 -4307 572
rect -4465 538 -4415 555
rect -4615 500 -4415 538
rect -4357 538 -4307 555
rect -4207 555 -4191 572
rect -4065 572 -3933 588
rect -4065 555 -4049 572
rect -4207 538 -4157 555
rect -4357 500 -4157 538
rect -4099 538 -4049 555
rect -3949 555 -3933 572
rect -3807 572 -3675 588
rect -3807 555 -3791 572
rect -3949 538 -3899 555
rect -4099 500 -3899 538
rect -3841 538 -3791 555
rect -3691 555 -3675 572
rect -3549 572 -3417 588
rect -3549 555 -3533 572
rect -3691 538 -3641 555
rect -3841 500 -3641 538
rect -3583 538 -3533 555
rect -3433 555 -3417 572
rect -3291 572 -3159 588
rect -3291 555 -3275 572
rect -3433 538 -3383 555
rect -3583 500 -3383 538
rect -3325 538 -3275 555
rect -3175 555 -3159 572
rect -3033 572 -2901 588
rect -3033 555 -3017 572
rect -3175 538 -3125 555
rect -3325 500 -3125 538
rect -3067 538 -3017 555
rect -2917 555 -2901 572
rect -2775 572 -2643 588
rect -2775 555 -2759 572
rect -2917 538 -2867 555
rect -3067 500 -2867 538
rect -2809 538 -2759 555
rect -2659 555 -2643 572
rect -2517 572 -2385 588
rect -2517 555 -2501 572
rect -2659 538 -2609 555
rect -2809 500 -2609 538
rect -2551 538 -2501 555
rect -2401 555 -2385 572
rect -2259 572 -2127 588
rect -2259 555 -2243 572
rect -2401 538 -2351 555
rect -2551 500 -2351 538
rect -2293 538 -2243 555
rect -2143 555 -2127 572
rect -2001 572 -1869 588
rect -2001 555 -1985 572
rect -2143 538 -2093 555
rect -2293 500 -2093 538
rect -2035 538 -1985 555
rect -1885 555 -1869 572
rect -1743 572 -1611 588
rect -1743 555 -1727 572
rect -1885 538 -1835 555
rect -2035 500 -1835 538
rect -1777 538 -1727 555
rect -1627 555 -1611 572
rect -1485 572 -1353 588
rect -1485 555 -1469 572
rect -1627 538 -1577 555
rect -1777 500 -1577 538
rect -1519 538 -1469 555
rect -1369 555 -1353 572
rect -1227 572 -1095 588
rect -1227 555 -1211 572
rect -1369 538 -1319 555
rect -1519 500 -1319 538
rect -1261 538 -1211 555
rect -1111 555 -1095 572
rect -969 572 -837 588
rect -969 555 -953 572
rect -1111 538 -1061 555
rect -1261 500 -1061 538
rect -1003 538 -953 555
rect -853 555 -837 572
rect -711 572 -579 588
rect -711 555 -695 572
rect -853 538 -803 555
rect -1003 500 -803 538
rect -745 538 -695 555
rect -595 555 -579 572
rect -453 572 -321 588
rect -453 555 -437 572
rect -595 538 -545 555
rect -745 500 -545 538
rect -487 538 -437 555
rect -337 555 -321 572
rect -195 572 -63 588
rect -195 555 -179 572
rect -337 538 -287 555
rect -487 500 -287 538
rect -229 538 -179 555
rect -79 555 -63 572
rect 63 572 195 588
rect 63 555 79 572
rect -79 538 -29 555
rect -229 500 -29 538
rect 29 538 79 555
rect 179 555 195 572
rect 321 572 453 588
rect 321 555 337 572
rect 179 538 229 555
rect 29 500 229 538
rect 287 538 337 555
rect 437 555 453 572
rect 579 572 711 588
rect 579 555 595 572
rect 437 538 487 555
rect 287 500 487 538
rect 545 538 595 555
rect 695 555 711 572
rect 837 572 969 588
rect 837 555 853 572
rect 695 538 745 555
rect 545 500 745 538
rect 803 538 853 555
rect 953 555 969 572
rect 1095 572 1227 588
rect 1095 555 1111 572
rect 953 538 1003 555
rect 803 500 1003 538
rect 1061 538 1111 555
rect 1211 555 1227 572
rect 1353 572 1485 588
rect 1353 555 1369 572
rect 1211 538 1261 555
rect 1061 500 1261 538
rect 1319 538 1369 555
rect 1469 555 1485 572
rect 1611 572 1743 588
rect 1611 555 1627 572
rect 1469 538 1519 555
rect 1319 500 1519 538
rect 1577 538 1627 555
rect 1727 555 1743 572
rect 1869 572 2001 588
rect 1869 555 1885 572
rect 1727 538 1777 555
rect 1577 500 1777 538
rect 1835 538 1885 555
rect 1985 555 2001 572
rect 2127 572 2259 588
rect 2127 555 2143 572
rect 1985 538 2035 555
rect 1835 500 2035 538
rect 2093 538 2143 555
rect 2243 555 2259 572
rect 2385 572 2517 588
rect 2385 555 2401 572
rect 2243 538 2293 555
rect 2093 500 2293 538
rect 2351 538 2401 555
rect 2501 555 2517 572
rect 2643 572 2775 588
rect 2643 555 2659 572
rect 2501 538 2551 555
rect 2351 500 2551 538
rect 2609 538 2659 555
rect 2759 555 2775 572
rect 2901 572 3033 588
rect 2901 555 2917 572
rect 2759 538 2809 555
rect 2609 500 2809 538
rect 2867 538 2917 555
rect 3017 555 3033 572
rect 3159 572 3291 588
rect 3159 555 3175 572
rect 3017 538 3067 555
rect 2867 500 3067 538
rect 3125 538 3175 555
rect 3275 555 3291 572
rect 3417 572 3549 588
rect 3417 555 3433 572
rect 3275 538 3325 555
rect 3125 500 3325 538
rect 3383 538 3433 555
rect 3533 555 3549 572
rect 3675 572 3807 588
rect 3675 555 3691 572
rect 3533 538 3583 555
rect 3383 500 3583 538
rect 3641 538 3691 555
rect 3791 555 3807 572
rect 3933 572 4065 588
rect 3933 555 3949 572
rect 3791 538 3841 555
rect 3641 500 3841 538
rect 3899 538 3949 555
rect 4049 555 4065 572
rect 4191 572 4323 588
rect 4191 555 4207 572
rect 4049 538 4099 555
rect 3899 500 4099 538
rect 4157 538 4207 555
rect 4307 555 4323 572
rect 4449 572 4581 588
rect 4449 555 4465 572
rect 4307 538 4357 555
rect 4157 500 4357 538
rect 4415 538 4465 555
rect 4565 555 4581 572
rect 4707 572 4839 588
rect 4707 555 4723 572
rect 4565 538 4615 555
rect 4415 500 4615 538
rect 4673 538 4723 555
rect 4823 555 4839 572
rect 4965 572 5097 588
rect 4965 555 4981 572
rect 4823 538 4873 555
rect 4673 500 4873 538
rect 4931 538 4981 555
rect 5081 555 5097 572
rect 5223 572 5355 588
rect 5223 555 5239 572
rect 5081 538 5131 555
rect 4931 500 5131 538
rect 5189 538 5239 555
rect 5339 555 5355 572
rect 5481 572 5613 588
rect 5481 555 5497 572
rect 5339 538 5389 555
rect 5189 500 5389 538
rect 5447 538 5497 555
rect 5597 555 5613 572
rect 5739 572 5871 588
rect 5739 555 5755 572
rect 5597 538 5647 555
rect 5447 500 5647 538
rect 5705 538 5755 555
rect 5855 555 5871 572
rect 5997 572 6129 588
rect 5997 555 6013 572
rect 5855 538 5905 555
rect 5705 500 5905 538
rect 5963 538 6013 555
rect 6113 555 6129 572
rect 6255 572 6387 588
rect 6255 555 6271 572
rect 6113 538 6163 555
rect 5963 500 6163 538
rect 6221 538 6271 555
rect 6371 555 6387 572
rect 6513 572 6645 588
rect 6513 555 6529 572
rect 6371 538 6421 555
rect 6221 500 6421 538
rect 6479 538 6529 555
rect 6629 555 6645 572
rect 6771 572 6903 588
rect 6771 555 6787 572
rect 6629 538 6679 555
rect 6479 500 6679 538
rect 6737 538 6787 555
rect 6887 555 6903 572
rect 6887 538 6937 555
rect 6737 500 6937 538
rect -6937 -538 -6737 -500
rect -6937 -555 -6887 -538
rect -6903 -572 -6887 -555
rect -6787 -555 -6737 -538
rect -6679 -538 -6479 -500
rect -6679 -555 -6629 -538
rect -6787 -572 -6771 -555
rect -6903 -588 -6771 -572
rect -6645 -572 -6629 -555
rect -6529 -555 -6479 -538
rect -6421 -538 -6221 -500
rect -6421 -555 -6371 -538
rect -6529 -572 -6513 -555
rect -6645 -588 -6513 -572
rect -6387 -572 -6371 -555
rect -6271 -555 -6221 -538
rect -6163 -538 -5963 -500
rect -6163 -555 -6113 -538
rect -6271 -572 -6255 -555
rect -6387 -588 -6255 -572
rect -6129 -572 -6113 -555
rect -6013 -555 -5963 -538
rect -5905 -538 -5705 -500
rect -5905 -555 -5855 -538
rect -6013 -572 -5997 -555
rect -6129 -588 -5997 -572
rect -5871 -572 -5855 -555
rect -5755 -555 -5705 -538
rect -5647 -538 -5447 -500
rect -5647 -555 -5597 -538
rect -5755 -572 -5739 -555
rect -5871 -588 -5739 -572
rect -5613 -572 -5597 -555
rect -5497 -555 -5447 -538
rect -5389 -538 -5189 -500
rect -5389 -555 -5339 -538
rect -5497 -572 -5481 -555
rect -5613 -588 -5481 -572
rect -5355 -572 -5339 -555
rect -5239 -555 -5189 -538
rect -5131 -538 -4931 -500
rect -5131 -555 -5081 -538
rect -5239 -572 -5223 -555
rect -5355 -588 -5223 -572
rect -5097 -572 -5081 -555
rect -4981 -555 -4931 -538
rect -4873 -538 -4673 -500
rect -4873 -555 -4823 -538
rect -4981 -572 -4965 -555
rect -5097 -588 -4965 -572
rect -4839 -572 -4823 -555
rect -4723 -555 -4673 -538
rect -4615 -538 -4415 -500
rect -4615 -555 -4565 -538
rect -4723 -572 -4707 -555
rect -4839 -588 -4707 -572
rect -4581 -572 -4565 -555
rect -4465 -555 -4415 -538
rect -4357 -538 -4157 -500
rect -4357 -555 -4307 -538
rect -4465 -572 -4449 -555
rect -4581 -588 -4449 -572
rect -4323 -572 -4307 -555
rect -4207 -555 -4157 -538
rect -4099 -538 -3899 -500
rect -4099 -555 -4049 -538
rect -4207 -572 -4191 -555
rect -4323 -588 -4191 -572
rect -4065 -572 -4049 -555
rect -3949 -555 -3899 -538
rect -3841 -538 -3641 -500
rect -3841 -555 -3791 -538
rect -3949 -572 -3933 -555
rect -4065 -588 -3933 -572
rect -3807 -572 -3791 -555
rect -3691 -555 -3641 -538
rect -3583 -538 -3383 -500
rect -3583 -555 -3533 -538
rect -3691 -572 -3675 -555
rect -3807 -588 -3675 -572
rect -3549 -572 -3533 -555
rect -3433 -555 -3383 -538
rect -3325 -538 -3125 -500
rect -3325 -555 -3275 -538
rect -3433 -572 -3417 -555
rect -3549 -588 -3417 -572
rect -3291 -572 -3275 -555
rect -3175 -555 -3125 -538
rect -3067 -538 -2867 -500
rect -3067 -555 -3017 -538
rect -3175 -572 -3159 -555
rect -3291 -588 -3159 -572
rect -3033 -572 -3017 -555
rect -2917 -555 -2867 -538
rect -2809 -538 -2609 -500
rect -2809 -555 -2759 -538
rect -2917 -572 -2901 -555
rect -3033 -588 -2901 -572
rect -2775 -572 -2759 -555
rect -2659 -555 -2609 -538
rect -2551 -538 -2351 -500
rect -2551 -555 -2501 -538
rect -2659 -572 -2643 -555
rect -2775 -588 -2643 -572
rect -2517 -572 -2501 -555
rect -2401 -555 -2351 -538
rect -2293 -538 -2093 -500
rect -2293 -555 -2243 -538
rect -2401 -572 -2385 -555
rect -2517 -588 -2385 -572
rect -2259 -572 -2243 -555
rect -2143 -555 -2093 -538
rect -2035 -538 -1835 -500
rect -2035 -555 -1985 -538
rect -2143 -572 -2127 -555
rect -2259 -588 -2127 -572
rect -2001 -572 -1985 -555
rect -1885 -555 -1835 -538
rect -1777 -538 -1577 -500
rect -1777 -555 -1727 -538
rect -1885 -572 -1869 -555
rect -2001 -588 -1869 -572
rect -1743 -572 -1727 -555
rect -1627 -555 -1577 -538
rect -1519 -538 -1319 -500
rect -1519 -555 -1469 -538
rect -1627 -572 -1611 -555
rect -1743 -588 -1611 -572
rect -1485 -572 -1469 -555
rect -1369 -555 -1319 -538
rect -1261 -538 -1061 -500
rect -1261 -555 -1211 -538
rect -1369 -572 -1353 -555
rect -1485 -588 -1353 -572
rect -1227 -572 -1211 -555
rect -1111 -555 -1061 -538
rect -1003 -538 -803 -500
rect -1003 -555 -953 -538
rect -1111 -572 -1095 -555
rect -1227 -588 -1095 -572
rect -969 -572 -953 -555
rect -853 -555 -803 -538
rect -745 -538 -545 -500
rect -745 -555 -695 -538
rect -853 -572 -837 -555
rect -969 -588 -837 -572
rect -711 -572 -695 -555
rect -595 -555 -545 -538
rect -487 -538 -287 -500
rect -487 -555 -437 -538
rect -595 -572 -579 -555
rect -711 -588 -579 -572
rect -453 -572 -437 -555
rect -337 -555 -287 -538
rect -229 -538 -29 -500
rect -229 -555 -179 -538
rect -337 -572 -321 -555
rect -453 -588 -321 -572
rect -195 -572 -179 -555
rect -79 -555 -29 -538
rect 29 -538 229 -500
rect 29 -555 79 -538
rect -79 -572 -63 -555
rect -195 -588 -63 -572
rect 63 -572 79 -555
rect 179 -555 229 -538
rect 287 -538 487 -500
rect 287 -555 337 -538
rect 179 -572 195 -555
rect 63 -588 195 -572
rect 321 -572 337 -555
rect 437 -555 487 -538
rect 545 -538 745 -500
rect 545 -555 595 -538
rect 437 -572 453 -555
rect 321 -588 453 -572
rect 579 -572 595 -555
rect 695 -555 745 -538
rect 803 -538 1003 -500
rect 803 -555 853 -538
rect 695 -572 711 -555
rect 579 -588 711 -572
rect 837 -572 853 -555
rect 953 -555 1003 -538
rect 1061 -538 1261 -500
rect 1061 -555 1111 -538
rect 953 -572 969 -555
rect 837 -588 969 -572
rect 1095 -572 1111 -555
rect 1211 -555 1261 -538
rect 1319 -538 1519 -500
rect 1319 -555 1369 -538
rect 1211 -572 1227 -555
rect 1095 -588 1227 -572
rect 1353 -572 1369 -555
rect 1469 -555 1519 -538
rect 1577 -538 1777 -500
rect 1577 -555 1627 -538
rect 1469 -572 1485 -555
rect 1353 -588 1485 -572
rect 1611 -572 1627 -555
rect 1727 -555 1777 -538
rect 1835 -538 2035 -500
rect 1835 -555 1885 -538
rect 1727 -572 1743 -555
rect 1611 -588 1743 -572
rect 1869 -572 1885 -555
rect 1985 -555 2035 -538
rect 2093 -538 2293 -500
rect 2093 -555 2143 -538
rect 1985 -572 2001 -555
rect 1869 -588 2001 -572
rect 2127 -572 2143 -555
rect 2243 -555 2293 -538
rect 2351 -538 2551 -500
rect 2351 -555 2401 -538
rect 2243 -572 2259 -555
rect 2127 -588 2259 -572
rect 2385 -572 2401 -555
rect 2501 -555 2551 -538
rect 2609 -538 2809 -500
rect 2609 -555 2659 -538
rect 2501 -572 2517 -555
rect 2385 -588 2517 -572
rect 2643 -572 2659 -555
rect 2759 -555 2809 -538
rect 2867 -538 3067 -500
rect 2867 -555 2917 -538
rect 2759 -572 2775 -555
rect 2643 -588 2775 -572
rect 2901 -572 2917 -555
rect 3017 -555 3067 -538
rect 3125 -538 3325 -500
rect 3125 -555 3175 -538
rect 3017 -572 3033 -555
rect 2901 -588 3033 -572
rect 3159 -572 3175 -555
rect 3275 -555 3325 -538
rect 3383 -538 3583 -500
rect 3383 -555 3433 -538
rect 3275 -572 3291 -555
rect 3159 -588 3291 -572
rect 3417 -572 3433 -555
rect 3533 -555 3583 -538
rect 3641 -538 3841 -500
rect 3641 -555 3691 -538
rect 3533 -572 3549 -555
rect 3417 -588 3549 -572
rect 3675 -572 3691 -555
rect 3791 -555 3841 -538
rect 3899 -538 4099 -500
rect 3899 -555 3949 -538
rect 3791 -572 3807 -555
rect 3675 -588 3807 -572
rect 3933 -572 3949 -555
rect 4049 -555 4099 -538
rect 4157 -538 4357 -500
rect 4157 -555 4207 -538
rect 4049 -572 4065 -555
rect 3933 -588 4065 -572
rect 4191 -572 4207 -555
rect 4307 -555 4357 -538
rect 4415 -538 4615 -500
rect 4415 -555 4465 -538
rect 4307 -572 4323 -555
rect 4191 -588 4323 -572
rect 4449 -572 4465 -555
rect 4565 -555 4615 -538
rect 4673 -538 4873 -500
rect 4673 -555 4723 -538
rect 4565 -572 4581 -555
rect 4449 -588 4581 -572
rect 4707 -572 4723 -555
rect 4823 -555 4873 -538
rect 4931 -538 5131 -500
rect 4931 -555 4981 -538
rect 4823 -572 4839 -555
rect 4707 -588 4839 -572
rect 4965 -572 4981 -555
rect 5081 -555 5131 -538
rect 5189 -538 5389 -500
rect 5189 -555 5239 -538
rect 5081 -572 5097 -555
rect 4965 -588 5097 -572
rect 5223 -572 5239 -555
rect 5339 -555 5389 -538
rect 5447 -538 5647 -500
rect 5447 -555 5497 -538
rect 5339 -572 5355 -555
rect 5223 -588 5355 -572
rect 5481 -572 5497 -555
rect 5597 -555 5647 -538
rect 5705 -538 5905 -500
rect 5705 -555 5755 -538
rect 5597 -572 5613 -555
rect 5481 -588 5613 -572
rect 5739 -572 5755 -555
rect 5855 -555 5905 -538
rect 5963 -538 6163 -500
rect 5963 -555 6013 -538
rect 5855 -572 5871 -555
rect 5739 -588 5871 -572
rect 5997 -572 6013 -555
rect 6113 -555 6163 -538
rect 6221 -538 6421 -500
rect 6221 -555 6271 -538
rect 6113 -572 6129 -555
rect 5997 -588 6129 -572
rect 6255 -572 6271 -555
rect 6371 -555 6421 -538
rect 6479 -538 6679 -500
rect 6479 -555 6529 -538
rect 6371 -572 6387 -555
rect 6255 -588 6387 -572
rect 6513 -572 6529 -555
rect 6629 -555 6679 -538
rect 6737 -538 6937 -500
rect 6737 -555 6787 -538
rect 6629 -572 6645 -555
rect 6513 -588 6645 -572
rect 6771 -572 6787 -555
rect 6887 -555 6937 -538
rect 6887 -572 6903 -555
rect 6771 -588 6903 -572
<< polycont >>
rect -6887 538 -6787 572
rect -6629 538 -6529 572
rect -6371 538 -6271 572
rect -6113 538 -6013 572
rect -5855 538 -5755 572
rect -5597 538 -5497 572
rect -5339 538 -5239 572
rect -5081 538 -4981 572
rect -4823 538 -4723 572
rect -4565 538 -4465 572
rect -4307 538 -4207 572
rect -4049 538 -3949 572
rect -3791 538 -3691 572
rect -3533 538 -3433 572
rect -3275 538 -3175 572
rect -3017 538 -2917 572
rect -2759 538 -2659 572
rect -2501 538 -2401 572
rect -2243 538 -2143 572
rect -1985 538 -1885 572
rect -1727 538 -1627 572
rect -1469 538 -1369 572
rect -1211 538 -1111 572
rect -953 538 -853 572
rect -695 538 -595 572
rect -437 538 -337 572
rect -179 538 -79 572
rect 79 538 179 572
rect 337 538 437 572
rect 595 538 695 572
rect 853 538 953 572
rect 1111 538 1211 572
rect 1369 538 1469 572
rect 1627 538 1727 572
rect 1885 538 1985 572
rect 2143 538 2243 572
rect 2401 538 2501 572
rect 2659 538 2759 572
rect 2917 538 3017 572
rect 3175 538 3275 572
rect 3433 538 3533 572
rect 3691 538 3791 572
rect 3949 538 4049 572
rect 4207 538 4307 572
rect 4465 538 4565 572
rect 4723 538 4823 572
rect 4981 538 5081 572
rect 5239 538 5339 572
rect 5497 538 5597 572
rect 5755 538 5855 572
rect 6013 538 6113 572
rect 6271 538 6371 572
rect 6529 538 6629 572
rect 6787 538 6887 572
rect -6887 -572 -6787 -538
rect -6629 -572 -6529 -538
rect -6371 -572 -6271 -538
rect -6113 -572 -6013 -538
rect -5855 -572 -5755 -538
rect -5597 -572 -5497 -538
rect -5339 -572 -5239 -538
rect -5081 -572 -4981 -538
rect -4823 -572 -4723 -538
rect -4565 -572 -4465 -538
rect -4307 -572 -4207 -538
rect -4049 -572 -3949 -538
rect -3791 -572 -3691 -538
rect -3533 -572 -3433 -538
rect -3275 -572 -3175 -538
rect -3017 -572 -2917 -538
rect -2759 -572 -2659 -538
rect -2501 -572 -2401 -538
rect -2243 -572 -2143 -538
rect -1985 -572 -1885 -538
rect -1727 -572 -1627 -538
rect -1469 -572 -1369 -538
rect -1211 -572 -1111 -538
rect -953 -572 -853 -538
rect -695 -572 -595 -538
rect -437 -572 -337 -538
rect -179 -572 -79 -538
rect 79 -572 179 -538
rect 337 -572 437 -538
rect 595 -572 695 -538
rect 853 -572 953 -538
rect 1111 -572 1211 -538
rect 1369 -572 1469 -538
rect 1627 -572 1727 -538
rect 1885 -572 1985 -538
rect 2143 -572 2243 -538
rect 2401 -572 2501 -538
rect 2659 -572 2759 -538
rect 2917 -572 3017 -538
rect 3175 -572 3275 -538
rect 3433 -572 3533 -538
rect 3691 -572 3791 -538
rect 3949 -572 4049 -538
rect 4207 -572 4307 -538
rect 4465 -572 4565 -538
rect 4723 -572 4823 -538
rect 4981 -572 5081 -538
rect 5239 -572 5339 -538
rect 5497 -572 5597 -538
rect 5755 -572 5855 -538
rect 6013 -572 6113 -538
rect 6271 -572 6371 -538
rect 6529 -572 6629 -538
rect 6787 -572 6887 -538
<< locali >>
rect -6903 538 -6887 572
rect -6787 538 -6771 572
rect -6645 538 -6629 572
rect -6529 538 -6513 572
rect -6387 538 -6371 572
rect -6271 538 -6255 572
rect -6129 538 -6113 572
rect -6013 538 -5997 572
rect -5871 538 -5855 572
rect -5755 538 -5739 572
rect -5613 538 -5597 572
rect -5497 538 -5481 572
rect -5355 538 -5339 572
rect -5239 538 -5223 572
rect -5097 538 -5081 572
rect -4981 538 -4965 572
rect -4839 538 -4823 572
rect -4723 538 -4707 572
rect -4581 538 -4565 572
rect -4465 538 -4449 572
rect -4323 538 -4307 572
rect -4207 538 -4191 572
rect -4065 538 -4049 572
rect -3949 538 -3933 572
rect -3807 538 -3791 572
rect -3691 538 -3675 572
rect -3549 538 -3533 572
rect -3433 538 -3417 572
rect -3291 538 -3275 572
rect -3175 538 -3159 572
rect -3033 538 -3017 572
rect -2917 538 -2901 572
rect -2775 538 -2759 572
rect -2659 538 -2643 572
rect -2517 538 -2501 572
rect -2401 538 -2385 572
rect -2259 538 -2243 572
rect -2143 538 -2127 572
rect -2001 538 -1985 572
rect -1885 538 -1869 572
rect -1743 538 -1727 572
rect -1627 538 -1611 572
rect -1485 538 -1469 572
rect -1369 538 -1353 572
rect -1227 538 -1211 572
rect -1111 538 -1095 572
rect -969 538 -953 572
rect -853 538 -837 572
rect -711 538 -695 572
rect -595 538 -579 572
rect -453 538 -437 572
rect -337 538 -321 572
rect -195 538 -179 572
rect -79 538 -63 572
rect 63 538 79 572
rect 179 538 195 572
rect 321 538 337 572
rect 437 538 453 572
rect 579 538 595 572
rect 695 538 711 572
rect 837 538 853 572
rect 953 538 969 572
rect 1095 538 1111 572
rect 1211 538 1227 572
rect 1353 538 1369 572
rect 1469 538 1485 572
rect 1611 538 1627 572
rect 1727 538 1743 572
rect 1869 538 1885 572
rect 1985 538 2001 572
rect 2127 538 2143 572
rect 2243 538 2259 572
rect 2385 538 2401 572
rect 2501 538 2517 572
rect 2643 538 2659 572
rect 2759 538 2775 572
rect 2901 538 2917 572
rect 3017 538 3033 572
rect 3159 538 3175 572
rect 3275 538 3291 572
rect 3417 538 3433 572
rect 3533 538 3549 572
rect 3675 538 3691 572
rect 3791 538 3807 572
rect 3933 538 3949 572
rect 4049 538 4065 572
rect 4191 538 4207 572
rect 4307 538 4323 572
rect 4449 538 4465 572
rect 4565 538 4581 572
rect 4707 538 4723 572
rect 4823 538 4839 572
rect 4965 538 4981 572
rect 5081 538 5097 572
rect 5223 538 5239 572
rect 5339 538 5355 572
rect 5481 538 5497 572
rect 5597 538 5613 572
rect 5739 538 5755 572
rect 5855 538 5871 572
rect 5997 538 6013 572
rect 6113 538 6129 572
rect 6255 538 6271 572
rect 6371 538 6387 572
rect 6513 538 6529 572
rect 6629 538 6645 572
rect 6771 538 6787 572
rect 6887 538 6903 572
rect -6983 488 -6949 504
rect -6983 -504 -6949 -488
rect -6725 488 -6691 504
rect -6725 -504 -6691 -488
rect -6467 488 -6433 504
rect -6467 -504 -6433 -488
rect -6209 488 -6175 504
rect -6209 -504 -6175 -488
rect -5951 488 -5917 504
rect -5951 -504 -5917 -488
rect -5693 488 -5659 504
rect -5693 -504 -5659 -488
rect -5435 488 -5401 504
rect -5435 -504 -5401 -488
rect -5177 488 -5143 504
rect -5177 -504 -5143 -488
rect -4919 488 -4885 504
rect -4919 -504 -4885 -488
rect -4661 488 -4627 504
rect -4661 -504 -4627 -488
rect -4403 488 -4369 504
rect -4403 -504 -4369 -488
rect -4145 488 -4111 504
rect -4145 -504 -4111 -488
rect -3887 488 -3853 504
rect -3887 -504 -3853 -488
rect -3629 488 -3595 504
rect -3629 -504 -3595 -488
rect -3371 488 -3337 504
rect -3371 -504 -3337 -488
rect -3113 488 -3079 504
rect -3113 -504 -3079 -488
rect -2855 488 -2821 504
rect -2855 -504 -2821 -488
rect -2597 488 -2563 504
rect -2597 -504 -2563 -488
rect -2339 488 -2305 504
rect -2339 -504 -2305 -488
rect -2081 488 -2047 504
rect -2081 -504 -2047 -488
rect -1823 488 -1789 504
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect 1789 488 1823 504
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -504 2081 -488
rect 2305 488 2339 504
rect 2305 -504 2339 -488
rect 2563 488 2597 504
rect 2563 -504 2597 -488
rect 2821 488 2855 504
rect 2821 -504 2855 -488
rect 3079 488 3113 504
rect 3079 -504 3113 -488
rect 3337 488 3371 504
rect 3337 -504 3371 -488
rect 3595 488 3629 504
rect 3595 -504 3629 -488
rect 3853 488 3887 504
rect 3853 -504 3887 -488
rect 4111 488 4145 504
rect 4111 -504 4145 -488
rect 4369 488 4403 504
rect 4369 -504 4403 -488
rect 4627 488 4661 504
rect 4627 -504 4661 -488
rect 4885 488 4919 504
rect 4885 -504 4919 -488
rect 5143 488 5177 504
rect 5143 -504 5177 -488
rect 5401 488 5435 504
rect 5401 -504 5435 -488
rect 5659 488 5693 504
rect 5659 -504 5693 -488
rect 5917 488 5951 504
rect 5917 -504 5951 -488
rect 6175 488 6209 504
rect 6175 -504 6209 -488
rect 6433 488 6467 504
rect 6433 -504 6467 -488
rect 6691 488 6725 504
rect 6691 -504 6725 -488
rect 6949 488 6983 504
rect 6949 -504 6983 -488
rect -6903 -572 -6887 -538
rect -6787 -572 -6771 -538
rect -6645 -572 -6629 -538
rect -6529 -572 -6513 -538
rect -6387 -572 -6371 -538
rect -6271 -572 -6255 -538
rect -6129 -572 -6113 -538
rect -6013 -572 -5997 -538
rect -5871 -572 -5855 -538
rect -5755 -572 -5739 -538
rect -5613 -572 -5597 -538
rect -5497 -572 -5481 -538
rect -5355 -572 -5339 -538
rect -5239 -572 -5223 -538
rect -5097 -572 -5081 -538
rect -4981 -572 -4965 -538
rect -4839 -572 -4823 -538
rect -4723 -572 -4707 -538
rect -4581 -572 -4565 -538
rect -4465 -572 -4449 -538
rect -4323 -572 -4307 -538
rect -4207 -572 -4191 -538
rect -4065 -572 -4049 -538
rect -3949 -572 -3933 -538
rect -3807 -572 -3791 -538
rect -3691 -572 -3675 -538
rect -3549 -572 -3533 -538
rect -3433 -572 -3417 -538
rect -3291 -572 -3275 -538
rect -3175 -572 -3159 -538
rect -3033 -572 -3017 -538
rect -2917 -572 -2901 -538
rect -2775 -572 -2759 -538
rect -2659 -572 -2643 -538
rect -2517 -572 -2501 -538
rect -2401 -572 -2385 -538
rect -2259 -572 -2243 -538
rect -2143 -572 -2127 -538
rect -2001 -572 -1985 -538
rect -1885 -572 -1869 -538
rect -1743 -572 -1727 -538
rect -1627 -572 -1611 -538
rect -1485 -572 -1469 -538
rect -1369 -572 -1353 -538
rect -1227 -572 -1211 -538
rect -1111 -572 -1095 -538
rect -969 -572 -953 -538
rect -853 -572 -837 -538
rect -711 -572 -695 -538
rect -595 -572 -579 -538
rect -453 -572 -437 -538
rect -337 -572 -321 -538
rect -195 -572 -179 -538
rect -79 -572 -63 -538
rect 63 -572 79 -538
rect 179 -572 195 -538
rect 321 -572 337 -538
rect 437 -572 453 -538
rect 579 -572 595 -538
rect 695 -572 711 -538
rect 837 -572 853 -538
rect 953 -572 969 -538
rect 1095 -572 1111 -538
rect 1211 -572 1227 -538
rect 1353 -572 1369 -538
rect 1469 -572 1485 -538
rect 1611 -572 1627 -538
rect 1727 -572 1743 -538
rect 1869 -572 1885 -538
rect 1985 -572 2001 -538
rect 2127 -572 2143 -538
rect 2243 -572 2259 -538
rect 2385 -572 2401 -538
rect 2501 -572 2517 -538
rect 2643 -572 2659 -538
rect 2759 -572 2775 -538
rect 2901 -572 2917 -538
rect 3017 -572 3033 -538
rect 3159 -572 3175 -538
rect 3275 -572 3291 -538
rect 3417 -572 3433 -538
rect 3533 -572 3549 -538
rect 3675 -572 3691 -538
rect 3791 -572 3807 -538
rect 3933 -572 3949 -538
rect 4049 -572 4065 -538
rect 4191 -572 4207 -538
rect 4307 -572 4323 -538
rect 4449 -572 4465 -538
rect 4565 -572 4581 -538
rect 4707 -572 4723 -538
rect 4823 -572 4839 -538
rect 4965 -572 4981 -538
rect 5081 -572 5097 -538
rect 5223 -572 5239 -538
rect 5339 -572 5355 -538
rect 5481 -572 5497 -538
rect 5597 -572 5613 -538
rect 5739 -572 5755 -538
rect 5855 -572 5871 -538
rect 5997 -572 6013 -538
rect 6113 -572 6129 -538
rect 6255 -572 6271 -538
rect 6371 -572 6387 -538
rect 6513 -572 6529 -538
rect 6629 -572 6645 -538
rect 6771 -572 6787 -538
rect 6887 -572 6903 -538
<< viali >>
rect -6871 538 -6803 572
rect -6613 538 -6545 572
rect -6355 538 -6287 572
rect -6097 538 -6029 572
rect -5839 538 -5771 572
rect -5581 538 -5513 572
rect -5323 538 -5255 572
rect -5065 538 -4997 572
rect -4807 538 -4739 572
rect -4549 538 -4481 572
rect -4291 538 -4223 572
rect -4033 538 -3965 572
rect -3775 538 -3707 572
rect -3517 538 -3449 572
rect -3259 538 -3191 572
rect -3001 538 -2933 572
rect -2743 538 -2675 572
rect -2485 538 -2417 572
rect -2227 538 -2159 572
rect -1969 538 -1901 572
rect -1711 538 -1643 572
rect -1453 538 -1385 572
rect -1195 538 -1127 572
rect -937 538 -869 572
rect -679 538 -611 572
rect -421 538 -353 572
rect -163 538 -95 572
rect 95 538 163 572
rect 353 538 421 572
rect 611 538 679 572
rect 869 538 937 572
rect 1127 538 1195 572
rect 1385 538 1453 572
rect 1643 538 1711 572
rect 1901 538 1969 572
rect 2159 538 2227 572
rect 2417 538 2485 572
rect 2675 538 2743 572
rect 2933 538 3001 572
rect 3191 538 3259 572
rect 3449 538 3517 572
rect 3707 538 3775 572
rect 3965 538 4033 572
rect 4223 538 4291 572
rect 4481 538 4549 572
rect 4739 538 4807 572
rect 4997 538 5065 572
rect 5255 538 5323 572
rect 5513 538 5581 572
rect 5771 538 5839 572
rect 6029 538 6097 572
rect 6287 538 6355 572
rect 6545 538 6613 572
rect 6803 538 6871 572
rect -6983 -488 -6949 488
rect -6725 -488 -6691 488
rect -6467 -488 -6433 488
rect -6209 -488 -6175 488
rect -5951 -488 -5917 488
rect -5693 -488 -5659 488
rect -5435 -488 -5401 488
rect -5177 -488 -5143 488
rect -4919 -488 -4885 488
rect -4661 -488 -4627 488
rect -4403 -488 -4369 488
rect -4145 -488 -4111 488
rect -3887 -488 -3853 488
rect -3629 -488 -3595 488
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect 3595 -488 3629 488
rect 3853 -488 3887 488
rect 4111 -488 4145 488
rect 4369 -488 4403 488
rect 4627 -488 4661 488
rect 4885 -488 4919 488
rect 5143 -488 5177 488
rect 5401 -488 5435 488
rect 5659 -488 5693 488
rect 5917 -488 5951 488
rect 6175 -488 6209 488
rect 6433 -488 6467 488
rect 6691 -488 6725 488
rect 6949 -488 6983 488
rect -6871 -572 -6803 -538
rect -6613 -572 -6545 -538
rect -6355 -572 -6287 -538
rect -6097 -572 -6029 -538
rect -5839 -572 -5771 -538
rect -5581 -572 -5513 -538
rect -5323 -572 -5255 -538
rect -5065 -572 -4997 -538
rect -4807 -572 -4739 -538
rect -4549 -572 -4481 -538
rect -4291 -572 -4223 -538
rect -4033 -572 -3965 -538
rect -3775 -572 -3707 -538
rect -3517 -572 -3449 -538
rect -3259 -572 -3191 -538
rect -3001 -572 -2933 -538
rect -2743 -572 -2675 -538
rect -2485 -572 -2417 -538
rect -2227 -572 -2159 -538
rect -1969 -572 -1901 -538
rect -1711 -572 -1643 -538
rect -1453 -572 -1385 -538
rect -1195 -572 -1127 -538
rect -937 -572 -869 -538
rect -679 -572 -611 -538
rect -421 -572 -353 -538
rect -163 -572 -95 -538
rect 95 -572 163 -538
rect 353 -572 421 -538
rect 611 -572 679 -538
rect 869 -572 937 -538
rect 1127 -572 1195 -538
rect 1385 -572 1453 -538
rect 1643 -572 1711 -538
rect 1901 -572 1969 -538
rect 2159 -572 2227 -538
rect 2417 -572 2485 -538
rect 2675 -572 2743 -538
rect 2933 -572 3001 -538
rect 3191 -572 3259 -538
rect 3449 -572 3517 -538
rect 3707 -572 3775 -538
rect 3965 -572 4033 -538
rect 4223 -572 4291 -538
rect 4481 -572 4549 -538
rect 4739 -572 4807 -538
rect 4997 -572 5065 -538
rect 5255 -572 5323 -538
rect 5513 -572 5581 -538
rect 5771 -572 5839 -538
rect 6029 -572 6097 -538
rect 6287 -572 6355 -538
rect 6545 -572 6613 -538
rect 6803 -572 6871 -538
<< metal1 >>
rect -6883 572 -6791 578
rect -6883 538 -6871 572
rect -6803 538 -6791 572
rect -6883 532 -6791 538
rect -6625 572 -6533 578
rect -6625 538 -6613 572
rect -6545 538 -6533 572
rect -6625 532 -6533 538
rect -6367 572 -6275 578
rect -6367 538 -6355 572
rect -6287 538 -6275 572
rect -6367 532 -6275 538
rect -6109 572 -6017 578
rect -6109 538 -6097 572
rect -6029 538 -6017 572
rect -6109 532 -6017 538
rect -5851 572 -5759 578
rect -5851 538 -5839 572
rect -5771 538 -5759 572
rect -5851 532 -5759 538
rect -5593 572 -5501 578
rect -5593 538 -5581 572
rect -5513 538 -5501 572
rect -5593 532 -5501 538
rect -5335 572 -5243 578
rect -5335 538 -5323 572
rect -5255 538 -5243 572
rect -5335 532 -5243 538
rect -5077 572 -4985 578
rect -5077 538 -5065 572
rect -4997 538 -4985 572
rect -5077 532 -4985 538
rect -4819 572 -4727 578
rect -4819 538 -4807 572
rect -4739 538 -4727 572
rect -4819 532 -4727 538
rect -4561 572 -4469 578
rect -4561 538 -4549 572
rect -4481 538 -4469 572
rect -4561 532 -4469 538
rect -4303 572 -4211 578
rect -4303 538 -4291 572
rect -4223 538 -4211 572
rect -4303 532 -4211 538
rect -4045 572 -3953 578
rect -4045 538 -4033 572
rect -3965 538 -3953 572
rect -4045 532 -3953 538
rect -3787 572 -3695 578
rect -3787 538 -3775 572
rect -3707 538 -3695 572
rect -3787 532 -3695 538
rect -3529 572 -3437 578
rect -3529 538 -3517 572
rect -3449 538 -3437 572
rect -3529 532 -3437 538
rect -3271 572 -3179 578
rect -3271 538 -3259 572
rect -3191 538 -3179 572
rect -3271 532 -3179 538
rect -3013 572 -2921 578
rect -3013 538 -3001 572
rect -2933 538 -2921 572
rect -3013 532 -2921 538
rect -2755 572 -2663 578
rect -2755 538 -2743 572
rect -2675 538 -2663 572
rect -2755 532 -2663 538
rect -2497 572 -2405 578
rect -2497 538 -2485 572
rect -2417 538 -2405 572
rect -2497 532 -2405 538
rect -2239 572 -2147 578
rect -2239 538 -2227 572
rect -2159 538 -2147 572
rect -2239 532 -2147 538
rect -1981 572 -1889 578
rect -1981 538 -1969 572
rect -1901 538 -1889 572
rect -1981 532 -1889 538
rect -1723 572 -1631 578
rect -1723 538 -1711 572
rect -1643 538 -1631 572
rect -1723 532 -1631 538
rect -1465 572 -1373 578
rect -1465 538 -1453 572
rect -1385 538 -1373 572
rect -1465 532 -1373 538
rect -1207 572 -1115 578
rect -1207 538 -1195 572
rect -1127 538 -1115 572
rect -1207 532 -1115 538
rect -949 572 -857 578
rect -949 538 -937 572
rect -869 538 -857 572
rect -949 532 -857 538
rect -691 572 -599 578
rect -691 538 -679 572
rect -611 538 -599 572
rect -691 532 -599 538
rect -433 572 -341 578
rect -433 538 -421 572
rect -353 538 -341 572
rect -433 532 -341 538
rect -175 572 -83 578
rect -175 538 -163 572
rect -95 538 -83 572
rect -175 532 -83 538
rect 83 572 175 578
rect 83 538 95 572
rect 163 538 175 572
rect 83 532 175 538
rect 341 572 433 578
rect 341 538 353 572
rect 421 538 433 572
rect 341 532 433 538
rect 599 572 691 578
rect 599 538 611 572
rect 679 538 691 572
rect 599 532 691 538
rect 857 572 949 578
rect 857 538 869 572
rect 937 538 949 572
rect 857 532 949 538
rect 1115 572 1207 578
rect 1115 538 1127 572
rect 1195 538 1207 572
rect 1115 532 1207 538
rect 1373 572 1465 578
rect 1373 538 1385 572
rect 1453 538 1465 572
rect 1373 532 1465 538
rect 1631 572 1723 578
rect 1631 538 1643 572
rect 1711 538 1723 572
rect 1631 532 1723 538
rect 1889 572 1981 578
rect 1889 538 1901 572
rect 1969 538 1981 572
rect 1889 532 1981 538
rect 2147 572 2239 578
rect 2147 538 2159 572
rect 2227 538 2239 572
rect 2147 532 2239 538
rect 2405 572 2497 578
rect 2405 538 2417 572
rect 2485 538 2497 572
rect 2405 532 2497 538
rect 2663 572 2755 578
rect 2663 538 2675 572
rect 2743 538 2755 572
rect 2663 532 2755 538
rect 2921 572 3013 578
rect 2921 538 2933 572
rect 3001 538 3013 572
rect 2921 532 3013 538
rect 3179 572 3271 578
rect 3179 538 3191 572
rect 3259 538 3271 572
rect 3179 532 3271 538
rect 3437 572 3529 578
rect 3437 538 3449 572
rect 3517 538 3529 572
rect 3437 532 3529 538
rect 3695 572 3787 578
rect 3695 538 3707 572
rect 3775 538 3787 572
rect 3695 532 3787 538
rect 3953 572 4045 578
rect 3953 538 3965 572
rect 4033 538 4045 572
rect 3953 532 4045 538
rect 4211 572 4303 578
rect 4211 538 4223 572
rect 4291 538 4303 572
rect 4211 532 4303 538
rect 4469 572 4561 578
rect 4469 538 4481 572
rect 4549 538 4561 572
rect 4469 532 4561 538
rect 4727 572 4819 578
rect 4727 538 4739 572
rect 4807 538 4819 572
rect 4727 532 4819 538
rect 4985 572 5077 578
rect 4985 538 4997 572
rect 5065 538 5077 572
rect 4985 532 5077 538
rect 5243 572 5335 578
rect 5243 538 5255 572
rect 5323 538 5335 572
rect 5243 532 5335 538
rect 5501 572 5593 578
rect 5501 538 5513 572
rect 5581 538 5593 572
rect 5501 532 5593 538
rect 5759 572 5851 578
rect 5759 538 5771 572
rect 5839 538 5851 572
rect 5759 532 5851 538
rect 6017 572 6109 578
rect 6017 538 6029 572
rect 6097 538 6109 572
rect 6017 532 6109 538
rect 6275 572 6367 578
rect 6275 538 6287 572
rect 6355 538 6367 572
rect 6275 532 6367 538
rect 6533 572 6625 578
rect 6533 538 6545 572
rect 6613 538 6625 572
rect 6533 532 6625 538
rect 6791 572 6883 578
rect 6791 538 6803 572
rect 6871 538 6883 572
rect 6791 532 6883 538
rect -6989 488 -6943 500
rect -6989 -488 -6983 488
rect -6949 -488 -6943 488
rect -6989 -500 -6943 -488
rect -6731 488 -6685 500
rect -6731 -488 -6725 488
rect -6691 -488 -6685 488
rect -6731 -500 -6685 -488
rect -6473 488 -6427 500
rect -6473 -488 -6467 488
rect -6433 -488 -6427 488
rect -6473 -500 -6427 -488
rect -6215 488 -6169 500
rect -6215 -488 -6209 488
rect -6175 -488 -6169 488
rect -6215 -500 -6169 -488
rect -5957 488 -5911 500
rect -5957 -488 -5951 488
rect -5917 -488 -5911 488
rect -5957 -500 -5911 -488
rect -5699 488 -5653 500
rect -5699 -488 -5693 488
rect -5659 -488 -5653 488
rect -5699 -500 -5653 -488
rect -5441 488 -5395 500
rect -5441 -488 -5435 488
rect -5401 -488 -5395 488
rect -5441 -500 -5395 -488
rect -5183 488 -5137 500
rect -5183 -488 -5177 488
rect -5143 -488 -5137 488
rect -5183 -500 -5137 -488
rect -4925 488 -4879 500
rect -4925 -488 -4919 488
rect -4885 -488 -4879 488
rect -4925 -500 -4879 -488
rect -4667 488 -4621 500
rect -4667 -488 -4661 488
rect -4627 -488 -4621 488
rect -4667 -500 -4621 -488
rect -4409 488 -4363 500
rect -4409 -488 -4403 488
rect -4369 -488 -4363 488
rect -4409 -500 -4363 -488
rect -4151 488 -4105 500
rect -4151 -488 -4145 488
rect -4111 -488 -4105 488
rect -4151 -500 -4105 -488
rect -3893 488 -3847 500
rect -3893 -488 -3887 488
rect -3853 -488 -3847 488
rect -3893 -500 -3847 -488
rect -3635 488 -3589 500
rect -3635 -488 -3629 488
rect -3595 -488 -3589 488
rect -3635 -500 -3589 -488
rect -3377 488 -3331 500
rect -3377 -488 -3371 488
rect -3337 -488 -3331 488
rect -3377 -500 -3331 -488
rect -3119 488 -3073 500
rect -3119 -488 -3113 488
rect -3079 -488 -3073 488
rect -3119 -500 -3073 -488
rect -2861 488 -2815 500
rect -2861 -488 -2855 488
rect -2821 -488 -2815 488
rect -2861 -500 -2815 -488
rect -2603 488 -2557 500
rect -2603 -488 -2597 488
rect -2563 -488 -2557 488
rect -2603 -500 -2557 -488
rect -2345 488 -2299 500
rect -2345 -488 -2339 488
rect -2305 -488 -2299 488
rect -2345 -500 -2299 -488
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
rect 2299 488 2345 500
rect 2299 -488 2305 488
rect 2339 -488 2345 488
rect 2299 -500 2345 -488
rect 2557 488 2603 500
rect 2557 -488 2563 488
rect 2597 -488 2603 488
rect 2557 -500 2603 -488
rect 2815 488 2861 500
rect 2815 -488 2821 488
rect 2855 -488 2861 488
rect 2815 -500 2861 -488
rect 3073 488 3119 500
rect 3073 -488 3079 488
rect 3113 -488 3119 488
rect 3073 -500 3119 -488
rect 3331 488 3377 500
rect 3331 -488 3337 488
rect 3371 -488 3377 488
rect 3331 -500 3377 -488
rect 3589 488 3635 500
rect 3589 -488 3595 488
rect 3629 -488 3635 488
rect 3589 -500 3635 -488
rect 3847 488 3893 500
rect 3847 -488 3853 488
rect 3887 -488 3893 488
rect 3847 -500 3893 -488
rect 4105 488 4151 500
rect 4105 -488 4111 488
rect 4145 -488 4151 488
rect 4105 -500 4151 -488
rect 4363 488 4409 500
rect 4363 -488 4369 488
rect 4403 -488 4409 488
rect 4363 -500 4409 -488
rect 4621 488 4667 500
rect 4621 -488 4627 488
rect 4661 -488 4667 488
rect 4621 -500 4667 -488
rect 4879 488 4925 500
rect 4879 -488 4885 488
rect 4919 -488 4925 488
rect 4879 -500 4925 -488
rect 5137 488 5183 500
rect 5137 -488 5143 488
rect 5177 -488 5183 488
rect 5137 -500 5183 -488
rect 5395 488 5441 500
rect 5395 -488 5401 488
rect 5435 -488 5441 488
rect 5395 -500 5441 -488
rect 5653 488 5699 500
rect 5653 -488 5659 488
rect 5693 -488 5699 488
rect 5653 -500 5699 -488
rect 5911 488 5957 500
rect 5911 -488 5917 488
rect 5951 -488 5957 488
rect 5911 -500 5957 -488
rect 6169 488 6215 500
rect 6169 -488 6175 488
rect 6209 -488 6215 488
rect 6169 -500 6215 -488
rect 6427 488 6473 500
rect 6427 -488 6433 488
rect 6467 -488 6473 488
rect 6427 -500 6473 -488
rect 6685 488 6731 500
rect 6685 -488 6691 488
rect 6725 -488 6731 488
rect 6685 -500 6731 -488
rect 6943 488 6989 500
rect 6943 -488 6949 488
rect 6983 -488 6989 488
rect 6943 -500 6989 -488
rect -6883 -538 -6791 -532
rect -6883 -572 -6871 -538
rect -6803 -572 -6791 -538
rect -6883 -578 -6791 -572
rect -6625 -538 -6533 -532
rect -6625 -572 -6613 -538
rect -6545 -572 -6533 -538
rect -6625 -578 -6533 -572
rect -6367 -538 -6275 -532
rect -6367 -572 -6355 -538
rect -6287 -572 -6275 -538
rect -6367 -578 -6275 -572
rect -6109 -538 -6017 -532
rect -6109 -572 -6097 -538
rect -6029 -572 -6017 -538
rect -6109 -578 -6017 -572
rect -5851 -538 -5759 -532
rect -5851 -572 -5839 -538
rect -5771 -572 -5759 -538
rect -5851 -578 -5759 -572
rect -5593 -538 -5501 -532
rect -5593 -572 -5581 -538
rect -5513 -572 -5501 -538
rect -5593 -578 -5501 -572
rect -5335 -538 -5243 -532
rect -5335 -572 -5323 -538
rect -5255 -572 -5243 -538
rect -5335 -578 -5243 -572
rect -5077 -538 -4985 -532
rect -5077 -572 -5065 -538
rect -4997 -572 -4985 -538
rect -5077 -578 -4985 -572
rect -4819 -538 -4727 -532
rect -4819 -572 -4807 -538
rect -4739 -572 -4727 -538
rect -4819 -578 -4727 -572
rect -4561 -538 -4469 -532
rect -4561 -572 -4549 -538
rect -4481 -572 -4469 -538
rect -4561 -578 -4469 -572
rect -4303 -538 -4211 -532
rect -4303 -572 -4291 -538
rect -4223 -572 -4211 -538
rect -4303 -578 -4211 -572
rect -4045 -538 -3953 -532
rect -4045 -572 -4033 -538
rect -3965 -572 -3953 -538
rect -4045 -578 -3953 -572
rect -3787 -538 -3695 -532
rect -3787 -572 -3775 -538
rect -3707 -572 -3695 -538
rect -3787 -578 -3695 -572
rect -3529 -538 -3437 -532
rect -3529 -572 -3517 -538
rect -3449 -572 -3437 -538
rect -3529 -578 -3437 -572
rect -3271 -538 -3179 -532
rect -3271 -572 -3259 -538
rect -3191 -572 -3179 -538
rect -3271 -578 -3179 -572
rect -3013 -538 -2921 -532
rect -3013 -572 -3001 -538
rect -2933 -572 -2921 -538
rect -3013 -578 -2921 -572
rect -2755 -538 -2663 -532
rect -2755 -572 -2743 -538
rect -2675 -572 -2663 -538
rect -2755 -578 -2663 -572
rect -2497 -538 -2405 -532
rect -2497 -572 -2485 -538
rect -2417 -572 -2405 -538
rect -2497 -578 -2405 -572
rect -2239 -538 -2147 -532
rect -2239 -572 -2227 -538
rect -2159 -572 -2147 -538
rect -2239 -578 -2147 -572
rect -1981 -538 -1889 -532
rect -1981 -572 -1969 -538
rect -1901 -572 -1889 -538
rect -1981 -578 -1889 -572
rect -1723 -538 -1631 -532
rect -1723 -572 -1711 -538
rect -1643 -572 -1631 -538
rect -1723 -578 -1631 -572
rect -1465 -538 -1373 -532
rect -1465 -572 -1453 -538
rect -1385 -572 -1373 -538
rect -1465 -578 -1373 -572
rect -1207 -538 -1115 -532
rect -1207 -572 -1195 -538
rect -1127 -572 -1115 -538
rect -1207 -578 -1115 -572
rect -949 -538 -857 -532
rect -949 -572 -937 -538
rect -869 -572 -857 -538
rect -949 -578 -857 -572
rect -691 -538 -599 -532
rect -691 -572 -679 -538
rect -611 -572 -599 -538
rect -691 -578 -599 -572
rect -433 -538 -341 -532
rect -433 -572 -421 -538
rect -353 -572 -341 -538
rect -433 -578 -341 -572
rect -175 -538 -83 -532
rect -175 -572 -163 -538
rect -95 -572 -83 -538
rect -175 -578 -83 -572
rect 83 -538 175 -532
rect 83 -572 95 -538
rect 163 -572 175 -538
rect 83 -578 175 -572
rect 341 -538 433 -532
rect 341 -572 353 -538
rect 421 -572 433 -538
rect 341 -578 433 -572
rect 599 -538 691 -532
rect 599 -572 611 -538
rect 679 -572 691 -538
rect 599 -578 691 -572
rect 857 -538 949 -532
rect 857 -572 869 -538
rect 937 -572 949 -538
rect 857 -578 949 -572
rect 1115 -538 1207 -532
rect 1115 -572 1127 -538
rect 1195 -572 1207 -538
rect 1115 -578 1207 -572
rect 1373 -538 1465 -532
rect 1373 -572 1385 -538
rect 1453 -572 1465 -538
rect 1373 -578 1465 -572
rect 1631 -538 1723 -532
rect 1631 -572 1643 -538
rect 1711 -572 1723 -538
rect 1631 -578 1723 -572
rect 1889 -538 1981 -532
rect 1889 -572 1901 -538
rect 1969 -572 1981 -538
rect 1889 -578 1981 -572
rect 2147 -538 2239 -532
rect 2147 -572 2159 -538
rect 2227 -572 2239 -538
rect 2147 -578 2239 -572
rect 2405 -538 2497 -532
rect 2405 -572 2417 -538
rect 2485 -572 2497 -538
rect 2405 -578 2497 -572
rect 2663 -538 2755 -532
rect 2663 -572 2675 -538
rect 2743 -572 2755 -538
rect 2663 -578 2755 -572
rect 2921 -538 3013 -532
rect 2921 -572 2933 -538
rect 3001 -572 3013 -538
rect 2921 -578 3013 -572
rect 3179 -538 3271 -532
rect 3179 -572 3191 -538
rect 3259 -572 3271 -538
rect 3179 -578 3271 -572
rect 3437 -538 3529 -532
rect 3437 -572 3449 -538
rect 3517 -572 3529 -538
rect 3437 -578 3529 -572
rect 3695 -538 3787 -532
rect 3695 -572 3707 -538
rect 3775 -572 3787 -538
rect 3695 -578 3787 -572
rect 3953 -538 4045 -532
rect 3953 -572 3965 -538
rect 4033 -572 4045 -538
rect 3953 -578 4045 -572
rect 4211 -538 4303 -532
rect 4211 -572 4223 -538
rect 4291 -572 4303 -538
rect 4211 -578 4303 -572
rect 4469 -538 4561 -532
rect 4469 -572 4481 -538
rect 4549 -572 4561 -538
rect 4469 -578 4561 -572
rect 4727 -538 4819 -532
rect 4727 -572 4739 -538
rect 4807 -572 4819 -538
rect 4727 -578 4819 -572
rect 4985 -538 5077 -532
rect 4985 -572 4997 -538
rect 5065 -572 5077 -538
rect 4985 -578 5077 -572
rect 5243 -538 5335 -532
rect 5243 -572 5255 -538
rect 5323 -572 5335 -538
rect 5243 -578 5335 -572
rect 5501 -538 5593 -532
rect 5501 -572 5513 -538
rect 5581 -572 5593 -538
rect 5501 -578 5593 -572
rect 5759 -538 5851 -532
rect 5759 -572 5771 -538
rect 5839 -572 5851 -538
rect 5759 -578 5851 -572
rect 6017 -538 6109 -532
rect 6017 -572 6029 -538
rect 6097 -572 6109 -538
rect 6017 -578 6109 -572
rect 6275 -538 6367 -532
rect 6275 -572 6287 -538
rect 6355 -572 6367 -538
rect 6275 -578 6367 -572
rect 6533 -538 6625 -532
rect 6533 -572 6545 -538
rect 6613 -572 6625 -538
rect 6533 -578 6625 -572
rect 6791 -538 6883 -532
rect 6791 -572 6803 -538
rect 6871 -572 6883 -538
rect 6791 -578 6883 -572
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 5 l 1 m 1 nf 54 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
