MACRO NMOS_S_54487678_X1_Y1
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN NMOS_S_54487678_X1_Y1 0 0 ;
  SIZE 2580 BY 7560 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 280 1460 560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260 4480 1460 4760 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 680 1860 6880 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 7225 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M2 ;
      RECT 690 700 1890 980 ;
    LAYER M2 ;
      RECT 690 6580 1890 6860 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6635 1375 6805 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V2 ;
      RECT 1645 765 1795 915 ;
    LAYER V2 ;
      RECT 1645 6645 1795 6795 ;
  END
END NMOS_S_54487678_X1_Y1
