magic
tech sky130A
magscale 1 2
timestamp 1624430562
<< nwell >>
rect -9000 40 9000 4500
<< pwell >>
rect -9000 -4500 9000 -40
<< mvpsubdiff >>
rect -8934 -118 8934 -106
rect -8934 -278 -8700 -118
rect 8700 -278 8934 -118
rect -8934 -290 8934 -278
rect -8934 -340 -8750 -290
rect -8934 -4200 -8922 -340
rect -8762 -4200 -8750 -340
rect -8934 -4250 -8750 -4200
rect 8750 -340 8934 -290
rect 8750 -4200 8762 -340
rect 8922 -4200 8934 -340
rect 8750 -4250 8934 -4200
rect -8934 -4262 8934 -4250
rect -8934 -4422 -8700 -4262
rect 8700 -4422 8934 -4262
rect -8934 -4434 8934 -4422
<< mvnsubdiff >>
rect -8934 4422 8934 4434
rect -8934 4262 -8700 4422
rect 8700 4262 8934 4422
rect -8934 4250 8934 4262
rect -8934 4200 -8750 4250
rect -8934 340 -8922 4200
rect -8762 340 -8750 4200
rect -8934 290 -8750 340
rect 8750 4200 8934 4250
rect 8750 340 8762 4200
rect 8922 340 8934 4200
rect 8750 290 8934 340
rect -8934 278 8934 290
rect -8934 118 -8700 278
rect 8700 118 8934 278
rect -8934 106 8934 118
<< mvpsubdiffcont >>
rect -8700 -278 8700 -118
rect -8922 -4200 -8762 -340
rect 8762 -4200 8922 -340
rect -8700 -4422 8700 -4262
<< mvnsubdiffcont >>
rect -8700 4262 8700 4422
rect -8922 340 -8762 4200
rect 8762 340 8922 4200
rect -8700 118 8700 278
<< locali >>
rect -8922 4200 -8762 4422
rect 8762 4200 8922 4422
rect -4839 3842 -1353 3868
rect -4839 3784 -2349 3842
rect -2291 3784 -1353 3842
rect -4839 3547 -1353 3784
rect -8922 118 -8762 340
rect 8762 118 8922 340
rect -8922 -340 -8762 -118
rect 8762 -340 8922 -118
rect -4323 -891 4323 -823
rect -4323 -949 -28 -891
rect 32 -949 4323 -891
rect -4323 -958 -27 -949
rect 29 -958 4323 -949
rect -4323 -992 4323 -958
rect -4323 -1028 -4191 -992
rect -3807 -1028 -3675 -992
rect -3291 -1028 -3159 -992
rect -3033 -1028 -2901 -992
rect -2775 -1028 -2643 -992
rect -2517 -1028 -2385 -992
rect -2259 -1028 -2127 -992
rect -2001 -1028 -1869 -992
rect -1227 -1028 -1095 -992
rect -969 -1028 -837 -992
rect -195 -1028 -63 -992
rect 63 -1028 195 -992
rect 837 -1028 969 -992
rect 1095 -1028 1227 -992
rect 1869 -1028 2001 -992
rect 2127 -1028 2259 -992
rect 2385 -1028 2517 -992
rect 2643 -1028 2775 -992
rect 2901 -1028 3033 -992
rect 3159 -1028 3291 -992
rect 3675 -1028 3807 -992
rect 4191 -1028 4323 -992
rect -1743 -2232 -1611 -2172
rect -1485 -2232 -1353 -2172
rect -711 -2232 -579 -2172
rect -453 -2232 -321 -2172
rect 321 -2232 453 -2172
rect 579 -2232 711 -2172
rect 1353 -2232 1485 -2172
rect 1611 -2232 1743 -2172
rect -1743 -2444 1743 -2232
rect -1743 -2502 255 -2444
rect 313 -2502 1743 -2444
rect -1743 -2511 1743 -2502
rect 236 -2512 336 -2511
rect -8922 -4422 -8762 -4200
rect 8762 -4422 8922 -4200
<< viali >>
rect -8762 4262 -8700 4422
rect -8700 4262 8700 4422
rect 8700 4262 8762 4422
rect -8922 477 -8762 4063
rect -2349 3784 -2291 3842
rect 8762 477 8922 4063
rect -8762 118 -8700 278
rect -8700 118 8700 278
rect 8700 118 8762 278
rect -8762 -278 -8700 -118
rect -8700 -278 8700 -118
rect 8700 -278 8762 -118
rect -8922 -4063 -8762 -477
rect -28 -949 32 -891
rect -27 -958 29 -949
rect 255 -2502 313 -2444
rect 8762 -4063 8922 -477
rect -8762 -4422 -8700 -4262
rect -8700 -4422 8700 -4262
rect 8700 -4422 8762 -4262
<< metal1 >>
rect -8928 4422 8928 4428
rect -8928 4262 -8762 4422
rect 8762 4262 8928 4422
rect -8928 4256 8928 4262
rect -8928 4063 -8756 4256
rect -8928 477 -8922 4063
rect -8762 477 -8756 4063
rect -8156 3956 -8146 4256
rect -5189 3587 -5131 4256
rect -4941 3600 -4931 3658
rect -4873 3600 -4863 3658
rect -5189 3541 -4985 3587
rect -5189 3500 -5131 3541
rect -4925 3500 -4879 3600
rect -4673 3500 -4615 4256
rect -4157 3500 -4099 4256
rect -3641 3500 -3583 4256
rect -3125 3500 -3067 4256
rect -2609 3500 -2551 4256
rect -2361 3842 -2279 3848
rect -2361 3784 -2349 3842
rect -2291 3784 -2279 3842
rect -2361 3778 -2279 3784
rect -2093 3500 -2035 4256
rect -1577 3500 -1519 4256
rect -1329 3600 -1319 3658
rect -1261 3600 -1251 3658
rect -1313 3500 -1267 3600
rect -1061 3587 -1003 4256
rect -1207 3541 -1003 3587
rect -1061 3500 -1003 3541
rect 2041 3587 2087 4256
rect 2299 3587 2345 4256
rect 2653 3947 2663 4007
rect 2755 3947 2765 4007
rect 2911 3947 2921 4007
rect 3013 3947 3023 4007
rect 2541 3620 2551 3678
rect 2609 3620 2619 3678
rect 2041 3541 2345 3587
rect 2041 3500 2087 3541
rect 2299 3500 2345 3541
rect 2557 3500 2603 3620
rect 2663 3587 2755 3947
rect 2921 3587 3013 3947
rect 3057 3620 3067 3678
rect 3125 3620 3135 3678
rect 3073 3500 3119 3620
rect 3331 3500 3377 4256
rect 3685 3947 3695 4007
rect 3787 3947 3797 4007
rect 3943 3947 3953 4007
rect 4045 3947 4055 4007
rect 3573 3788 3583 3846
rect 3641 3788 3651 3846
rect 3589 3500 3635 3788
rect 3695 3587 3787 3947
rect 3953 3587 4045 3947
rect 4089 3788 4099 3846
rect 4157 3788 4167 3846
rect 4105 3500 4151 3788
rect 4363 3500 4409 4256
rect 4717 3947 4727 4007
rect 4819 3947 4829 4007
rect 4975 3947 4985 4007
rect 5077 3947 5087 4007
rect 4605 3620 4615 3678
rect 4673 3620 4683 3678
rect 4621 3500 4667 3620
rect 4727 3587 4819 3947
rect 4985 3587 5077 3947
rect 5121 3620 5131 3678
rect 5189 3620 5199 3678
rect 5137 3500 5183 3620
rect 5395 3500 5441 4256
rect 5749 3947 5759 4007
rect 5851 3947 5861 4007
rect 6007 3947 6017 4007
rect 6109 3947 6119 4007
rect 5638 3788 5648 3846
rect 5706 3788 5716 3846
rect 5653 3500 5699 3788
rect 5759 3587 5851 3947
rect 6017 3587 6109 3947
rect 6153 3788 6163 3846
rect 6221 3788 6231 3846
rect 6169 3500 6215 3788
rect 6427 3587 6473 4256
rect 6685 3587 6731 4256
rect 8146 3956 8156 4256
rect 8756 4063 8928 4256
rect 6427 3541 6731 3587
rect 6427 3500 6473 3541
rect 6685 3500 6731 3541
rect -4409 2373 -4363 2500
rect -3893 2373 -3847 2500
rect -3377 2373 -3331 2500
rect -2861 2373 -2815 2500
rect -2345 2373 -2299 2500
rect -1829 2373 -1783 2500
rect 2815 2435 2861 2500
rect -4409 2257 63 2373
rect 2405 2317 2497 2413
rect 2799 2377 2809 2435
rect 2867 2377 2877 2435
rect 3179 2317 3271 2413
rect 3437 2317 3529 2413
rect 3847 2317 3893 2500
rect 4879 2435 4925 2500
rect 4211 2317 4303 2413
rect 4469 2317 4561 2413
rect 4863 2377 4873 2435
rect 4931 2377 4941 2435
rect 5243 2317 5335 2413
rect 5501 2317 5593 2413
rect 5911 2317 5957 2500
rect 6275 2317 6367 2413
rect 2405 2257 7194 2317
rect -63 2217 63 2257
rect 7114 2239 7194 2257
rect -6989 2137 6989 2217
rect 7114 2181 7125 2239
rect 7183 2181 7194 2239
rect -6989 1887 -6943 2137
rect -6731 1887 -6685 2137
rect -6635 1917 -6625 1977
rect -6533 1917 -6523 1977
rect -6377 1917 -6367 1977
rect -6275 1917 -6265 1977
rect -6625 1887 -6533 1917
rect -6367 1887 -6275 1917
rect -6989 1842 -6685 1887
rect -6989 1800 -6943 1842
rect -6731 1800 -6685 1842
rect -6215 1800 -6169 2137
rect -6119 2037 -6109 2097
rect -6017 2037 -6007 2097
rect -5861 2037 -5851 2097
rect -5759 2037 -5749 2097
rect -6109 1887 -6017 2037
rect -5851 1887 -5759 2037
rect -5699 1800 -5653 2137
rect -5603 1917 -5593 1977
rect -5501 1917 -5491 1977
rect -5345 1917 -5335 1977
rect -5243 1917 -5233 1977
rect -5593 1887 -5501 1917
rect -5335 1887 -5243 1917
rect -5183 1800 -5137 2137
rect -5087 2037 -5077 2097
rect -4985 2037 -4975 2097
rect -4829 2037 -4819 2097
rect -4727 2037 -4717 2097
rect -5077 1887 -4985 2037
rect -4819 1887 -4727 2037
rect -4667 1800 -4621 2137
rect -4571 1917 -4561 1977
rect -4469 1917 -4459 1977
rect -4313 1917 -4303 1977
rect -4211 1917 -4201 1977
rect -4561 1887 -4469 1917
rect -4303 1887 -4211 1917
rect -4151 1800 -4105 2137
rect -4055 2037 -4045 2097
rect -3953 2037 -3943 2097
rect -3797 2037 -3787 2097
rect -3695 2037 -3685 2097
rect -4045 1887 -3953 2037
rect -3787 1887 -3695 2037
rect -3635 1800 -3589 2137
rect -3539 1917 -3529 1977
rect -3437 1917 -3427 1977
rect -3281 1917 -3271 1977
rect -3179 1917 -3169 1977
rect -3529 1887 -3437 1917
rect -3271 1887 -3179 1917
rect -3119 1800 -3073 2137
rect -3023 2037 -3013 2097
rect -2921 2037 -2911 2097
rect -2765 2037 -2755 2097
rect -2663 2037 -2653 2097
rect -3013 1887 -2921 2037
rect -2755 1887 -2663 2037
rect -2603 1800 -2557 2137
rect -2507 1917 -2497 1977
rect -2405 1917 -2395 1977
rect -2249 1917 -2239 1977
rect -2147 1917 -2137 1977
rect -2497 1887 -2405 1917
rect -2239 1887 -2147 1917
rect -2087 1800 -2041 2137
rect -1991 2037 -1981 2097
rect -1889 2037 -1879 2097
rect -1733 2037 -1723 2097
rect -1631 2037 -1621 2097
rect -1981 1887 -1889 2037
rect -1723 1887 -1631 2037
rect -1571 1800 -1525 2137
rect -1475 1917 -1465 1977
rect -1373 1917 -1363 1977
rect -1217 1917 -1207 1977
rect -1115 1917 -1105 1977
rect -1465 1887 -1373 1917
rect -1207 1887 -1115 1917
rect -1055 1800 -1009 2137
rect -959 2037 -949 2097
rect -857 2037 -847 2097
rect -701 2037 -691 2097
rect -599 2037 -589 2097
rect -949 1887 -857 2037
rect -691 1887 -599 2037
rect -539 1800 -493 2137
rect 331 2037 341 2097
rect 433 2037 443 2097
rect -443 1917 -433 1977
rect -341 1917 -331 1977
rect -433 1887 -341 1917
rect 341 1887 433 2037
rect 493 1800 539 2137
rect 589 1917 599 1977
rect 691 1917 701 1977
rect 847 1917 857 1977
rect 949 1917 959 1977
rect 599 1887 691 1917
rect 857 1887 949 1917
rect 1009 1800 1055 2137
rect 1105 2037 1115 2097
rect 1207 2037 1217 2097
rect 1363 2037 1373 2097
rect 1465 2037 1475 2097
rect 1115 1887 1207 2037
rect 1373 1887 1465 2037
rect 1525 1800 1571 2137
rect 1621 1917 1631 1977
rect 1723 1917 1733 1977
rect 1879 1917 1889 1977
rect 1981 1917 1991 1977
rect 1631 1887 1723 1917
rect 1889 1887 1981 1917
rect 2041 1800 2087 2137
rect 2137 2037 2147 2097
rect 2239 2037 2249 2097
rect 2395 2037 2405 2097
rect 2497 2037 2507 2097
rect 2147 1887 2239 2037
rect 2405 1887 2497 2037
rect 2557 1800 2603 2137
rect 2653 1917 2663 1977
rect 2755 1917 2765 1977
rect 2911 1917 2921 1977
rect 3013 1917 3023 1977
rect 2663 1887 2755 1917
rect 2921 1887 3013 1917
rect 3073 1800 3119 2137
rect 3169 2037 3179 2097
rect 3271 2037 3281 2097
rect 3427 2037 3437 2097
rect 3529 2037 3539 2097
rect 3179 1887 3271 2037
rect 3437 1887 3529 2037
rect 3589 1800 3635 2137
rect 3685 1917 3695 1977
rect 3787 1917 3797 1977
rect 3943 1917 3953 1977
rect 4045 1917 4055 1977
rect 3695 1887 3787 1917
rect 3953 1887 4045 1917
rect 4105 1800 4151 2137
rect 4201 2037 4211 2097
rect 4303 2037 4313 2097
rect 4459 2037 4469 2097
rect 4561 2037 4571 2097
rect 4211 1887 4303 2037
rect 4469 1887 4561 2037
rect 4621 1800 4667 2137
rect 4717 1917 4727 1977
rect 4819 1917 4829 1977
rect 4975 1917 4985 1977
rect 5077 1917 5087 1977
rect 4727 1887 4819 1917
rect 4985 1887 5077 1917
rect 5137 1800 5183 2137
rect 5233 2037 5243 2097
rect 5335 2037 5345 2097
rect 5491 2037 5501 2097
rect 5593 2037 5603 2097
rect 5243 1887 5335 2037
rect 5501 1887 5593 2037
rect 5653 1800 5699 2137
rect 5749 1917 5759 1977
rect 5851 1917 5861 1977
rect 6007 1917 6017 1977
rect 6109 1917 6119 1977
rect 5759 1887 5851 1917
rect 6017 1887 6109 1917
rect 6169 1800 6215 2137
rect 6265 2037 6275 2097
rect 6367 2037 6377 2097
rect 6523 2037 6533 2097
rect 6625 2037 6635 2097
rect 6275 1887 6367 2037
rect 6533 1887 6625 2037
rect 6685 1886 6731 2137
rect 6943 1886 6989 2137
rect 6685 1841 6989 1886
rect 6685 1800 6731 1841
rect 6943 1800 6989 1841
rect -6473 560 -6427 800
rect -5957 700 -5911 800
rect -5973 642 -5963 700
rect -5905 642 -5895 700
rect -5441 560 -5395 800
rect -4925 700 -4879 800
rect -4941 642 -4931 700
rect -4873 642 -4863 700
rect -4409 560 -4363 800
rect -3893 700 -3847 800
rect -3909 642 -3899 700
rect -3841 642 -3831 700
rect -3377 561 -3331 801
rect -2861 700 -2815 800
rect -2877 642 -2867 700
rect -2809 642 -2799 700
rect -6489 502 -6479 560
rect -6421 502 -6411 560
rect -5457 502 -5447 560
rect -5389 502 -5379 560
rect -4425 502 -4415 560
rect -4357 502 -4347 560
rect -3393 503 -3383 561
rect -3325 503 -3315 561
rect -2345 560 -2299 800
rect -1829 700 -1783 800
rect -1845 642 -1835 700
rect -1777 642 -1767 700
rect -1313 560 -1267 800
rect -797 700 -751 800
rect -813 642 -803 700
rect -745 642 -735 700
rect -281 560 -235 800
rect -23 759 23 800
rect -175 713 175 759
rect -2361 502 -2351 560
rect -2293 502 -2283 560
rect -1329 502 -1319 560
rect -1261 502 -1251 560
rect -297 502 -287 560
rect -229 502 -219 560
rect -8928 284 -8756 477
rect -23 401 23 713
rect 235 700 281 800
rect 219 642 229 700
rect 287 642 297 700
rect 219 401 297 642
rect 751 561 797 801
rect 1267 700 1313 800
rect 1251 642 1261 700
rect 1319 642 1329 700
rect 735 503 745 561
rect 803 503 813 561
rect 1783 560 1829 800
rect 2299 700 2345 800
rect 2283 642 2293 700
rect 2351 642 2361 700
rect 2815 560 2861 800
rect 3331 700 3377 800
rect 3315 642 3325 700
rect 3383 642 3393 700
rect 3847 560 3893 800
rect 4363 700 4409 800
rect 4347 642 4357 700
rect 4415 642 4425 700
rect 4879 560 4925 800
rect 5395 700 5441 800
rect 5379 642 5389 700
rect 5447 642 5457 700
rect 5911 560 5957 800
rect 6427 700 6473 800
rect 6411 642 6421 700
rect 6479 642 6489 700
rect 1767 502 1777 560
rect 1835 502 1845 560
rect 2799 502 2809 560
rect 2867 502 2877 560
rect 3831 502 3841 560
rect 3899 502 3909 560
rect 4863 502 4873 560
rect 4931 502 4941 560
rect 5895 502 5905 560
rect 5963 502 5973 560
rect -39 343 -29 401
rect 29 343 39 401
rect 219 343 229 401
rect 287 343 297 401
rect 8756 477 8762 4063
rect 8922 477 8928 4063
rect 8756 284 8928 477
rect -8928 278 8928 284
rect -8928 118 -8762 278
rect 8762 118 8928 278
rect -8928 112 8928 118
rect -8928 -118 8928 -112
rect -8928 -278 -8762 -118
rect 8762 -278 8928 -118
rect -8928 -284 8928 -278
rect -8928 -477 -8756 -284
rect -8928 -4063 -8922 -477
rect -8762 -4063 -8756 -477
rect -298 -378 -287 -320
rect -229 -378 -218 -320
rect -1587 -646 -1577 -588
rect -1519 -646 -1509 -588
rect -3909 -764 -3899 -706
rect -3841 -764 -3831 -706
rect -2877 -764 -2867 -706
rect -2809 -764 -2799 -706
rect -1845 -764 -1835 -706
rect -1777 -764 -1767 -706
rect -3893 -1100 -3847 -764
rect -3393 -1000 -3383 -942
rect -3325 -1000 -3315 -942
rect -3377 -1100 -3331 -1000
rect -2861 -1100 -2815 -764
rect -2361 -1000 -2351 -942
rect -2293 -1000 -2283 -942
rect -2345 -1100 -2299 -1000
rect -1829 -1100 -1783 -764
rect -1571 -1100 -1525 -646
rect -1329 -764 -1319 -706
rect -1261 -764 -1251 -706
rect -1313 -1100 -1267 -764
rect -555 -882 -545 -824
rect -487 -882 -477 -824
rect -813 -1000 -803 -942
rect -745 -1000 -735 -942
rect -797 -1100 -751 -1000
rect -539 -1100 -493 -882
rect -298 -942 -218 -378
rect -298 -1000 -287 -942
rect -229 -1000 -218 -942
rect -40 -378 -29 -320
rect 29 -378 40 -320
rect -40 -891 40 -378
rect 218 -378 229 -320
rect 287 -378 297 -320
rect 218 -460 297 -378
rect 218 -706 298 -460
rect 8756 -477 8928 -284
rect 605 -588 685 -578
rect 477 -646 487 -588
rect 545 -646 555 -588
rect 605 -646 616 -588
rect 674 -646 685 -588
rect 218 -764 229 -706
rect 287 -764 298 -706
rect -40 -949 -28 -891
rect 32 -949 40 -891
rect -40 -958 -27 -949
rect 29 -958 40 -949
rect -40 -967 40 -958
rect -33 -970 35 -967
rect -281 -1100 -235 -1000
rect 235 -1100 281 -764
rect 493 -1100 539 -646
rect 605 -825 685 -646
rect 735 -764 745 -706
rect 803 -764 813 -706
rect 2283 -764 2293 -706
rect 2351 -764 2361 -706
rect 3315 -764 3325 -706
rect 3383 -764 3393 -706
rect 605 -883 616 -825
rect 674 -883 685 -825
rect 751 -1100 797 -764
rect 1509 -882 1519 -824
rect 1577 -882 1587 -824
rect 1251 -1000 1261 -942
rect 1319 -1000 1329 -942
rect 1267 -1100 1313 -1000
rect 1525 -1100 1571 -882
rect 1767 -1000 1777 -942
rect 1835 -1000 1845 -942
rect 1783 -1100 1829 -1000
rect 2299 -1100 2345 -764
rect 2799 -1000 2809 -942
rect 2867 -1000 2877 -942
rect 2815 -1100 2861 -1000
rect 3331 -1100 3377 -764
rect 3831 -1000 3841 -942
rect 3899 -1000 3909 -942
rect 3847 -1100 3893 -1000
rect -4667 -2228 -4621 -2100
rect -4409 -2130 -4363 -2100
rect -4561 -2228 -4469 -2178
rect -4425 -2188 -4415 -2130
rect -4357 -2188 -4211 -2130
rect -4151 -2228 -4105 -2100
rect -4045 -2228 -3953 -2178
rect -3635 -2228 -3589 -2100
rect -3529 -2228 -3437 -2178
rect -3119 -2228 -3073 -2100
rect -2603 -2228 -2557 -2100
rect -2087 -2228 -2041 -2100
rect -1055 -2228 -1009 -2100
rect -23 -2228 23 -2100
rect 1009 -2228 1055 -2100
rect 2041 -2228 2087 -2100
rect 2557 -2228 2603 -2100
rect 3073 -2228 3119 -2100
rect 3437 -2228 3529 -2178
rect 3589 -2228 3635 -2100
rect 3953 -2228 4045 -2178
rect 4105 -2228 4151 -2100
rect 4363 -2130 4409 -2100
rect 4211 -2188 4357 -2130
rect 4415 -2188 4425 -2130
rect 4469 -2228 4561 -2178
rect 4621 -2228 4667 -2100
rect -4667 -2328 4667 -2228
rect -8928 -4256 -8756 -4063
rect -8156 -4256 -8146 -3956
rect -4667 -4256 -4567 -2328
rect -2372 -4256 -2272 -2328
rect -50 -4256 50 -2328
rect 243 -2444 325 -2438
rect 243 -2502 255 -2444
rect 313 -2502 325 -2444
rect 243 -2508 325 -2502
rect 2272 -4256 2372 -2328
rect 4567 -4256 4667 -2328
rect 8146 -4256 8156 -3956
rect 8756 -4063 8762 -477
rect 8922 -4063 8928 -477
rect 8756 -4256 8928 -4063
rect -8928 -4262 8928 -4256
rect -8928 -4422 -8762 -4262
rect 8762 -4422 8928 -4262
rect -8928 -4428 8928 -4422
<< via1 >>
rect -8756 3956 -8156 4256
rect -4931 3600 -4873 3658
rect -2349 3784 -2291 3842
rect -1319 3600 -1261 3658
rect 2663 3947 2755 4007
rect 2921 3947 3013 4007
rect 2551 3620 2609 3678
rect 3067 3620 3125 3678
rect 3695 3947 3787 4007
rect 3953 3947 4045 4007
rect 3583 3788 3641 3846
rect 4099 3788 4157 3846
rect 4727 3947 4819 4007
rect 4985 3947 5077 4007
rect 4615 3620 4673 3678
rect 5131 3620 5189 3678
rect 5759 3947 5851 4007
rect 6017 3947 6109 4007
rect 5648 3788 5706 3846
rect 6163 3788 6221 3846
rect 8156 3956 8756 4256
rect 2809 2377 2867 2435
rect 4873 2377 4931 2435
rect 7125 2181 7183 2239
rect -6625 1917 -6533 1977
rect -6367 1917 -6275 1977
rect -6109 2037 -6017 2097
rect -5851 2037 -5759 2097
rect -5593 1917 -5501 1977
rect -5335 1917 -5243 1977
rect -5077 2037 -4985 2097
rect -4819 2037 -4727 2097
rect -4561 1917 -4469 1977
rect -4303 1917 -4211 1977
rect -4045 2037 -3953 2097
rect -3787 2037 -3695 2097
rect -3529 1917 -3437 1977
rect -3271 1917 -3179 1977
rect -3013 2037 -2921 2097
rect -2755 2037 -2663 2097
rect -2497 1917 -2405 1977
rect -2239 1917 -2147 1977
rect -1981 2037 -1889 2097
rect -1723 2037 -1631 2097
rect -1465 1917 -1373 1977
rect -1207 1917 -1115 1977
rect -949 2037 -857 2097
rect -691 2037 -599 2097
rect 341 2037 433 2097
rect -433 1917 -341 1977
rect 599 1917 691 1977
rect 857 1917 949 1977
rect 1115 2037 1207 2097
rect 1373 2037 1465 2097
rect 1631 1917 1723 1977
rect 1889 1917 1981 1977
rect 2147 2037 2239 2097
rect 2405 2037 2497 2097
rect 2663 1917 2755 1977
rect 2921 1917 3013 1977
rect 3179 2037 3271 2097
rect 3437 2037 3529 2097
rect 3695 1917 3787 1977
rect 3953 1917 4045 1977
rect 4211 2037 4303 2097
rect 4469 2037 4561 2097
rect 4727 1917 4819 1977
rect 4985 1917 5077 1977
rect 5243 2037 5335 2097
rect 5501 2037 5593 2097
rect 5759 1917 5851 1977
rect 6017 1917 6109 1977
rect 6275 2037 6367 2097
rect 6533 2037 6625 2097
rect -5963 642 -5905 700
rect -4931 642 -4873 700
rect -3899 642 -3841 700
rect -2867 642 -2809 700
rect -6479 502 -6421 560
rect -5447 502 -5389 560
rect -4415 502 -4357 560
rect -3383 503 -3325 561
rect -1835 642 -1777 700
rect -803 642 -745 700
rect -2351 502 -2293 560
rect -1319 502 -1261 560
rect -287 502 -229 560
rect 229 642 287 700
rect 1261 642 1319 700
rect 745 503 803 561
rect 2293 642 2351 700
rect 3325 642 3383 700
rect 4357 642 4415 700
rect 5389 642 5447 700
rect 6421 642 6479 700
rect 1777 502 1835 560
rect 2809 502 2867 560
rect 3841 502 3899 560
rect 4873 502 4931 560
rect 5905 502 5963 560
rect -29 343 29 401
rect 229 343 287 401
rect -287 -378 -229 -320
rect -1577 -646 -1519 -588
rect -3899 -764 -3841 -706
rect -2867 -764 -2809 -706
rect -1835 -764 -1777 -706
rect -3383 -1000 -3325 -942
rect -2351 -1000 -2293 -942
rect -1319 -764 -1261 -706
rect -545 -882 -487 -824
rect -803 -1000 -745 -942
rect -287 -1000 -229 -942
rect -29 -378 29 -320
rect 229 -378 287 -320
rect 487 -646 545 -588
rect 616 -646 674 -588
rect 229 -764 287 -706
rect 745 -764 803 -706
rect 2293 -764 2351 -706
rect 3325 -764 3383 -706
rect 616 -883 674 -825
rect 1519 -882 1577 -824
rect 1261 -1000 1319 -942
rect 1777 -1000 1835 -942
rect 2809 -1000 2867 -942
rect 3841 -1000 3899 -942
rect -4415 -2188 -4357 -2130
rect 4357 -2188 4415 -2130
rect -8756 -4256 -8156 -3956
rect 255 -2502 313 -2444
rect 8156 -4256 8756 -3956
<< metal2 >>
rect -8756 4256 -8156 4266
rect 8156 4256 8756 4266
rect -8756 3946 -8156 3956
rect 2663 4007 6384 4017
rect 2755 3947 2921 4007
rect 3013 3947 3695 4007
rect 3787 3947 3953 4007
rect 4045 3947 4727 4007
rect 4819 3947 4985 4007
rect 5077 3947 5759 4007
rect 5851 3947 6017 4007
rect 6109 3947 6384 4007
rect 2663 3937 6384 3947
rect 8156 3946 8756 3956
rect -2349 3842 -2291 3852
rect -7756 3708 -3033 3828
rect -2349 3774 -2291 3784
rect 3583 3846 6221 3856
rect 3641 3796 4099 3846
rect 3583 3778 3641 3788
rect 4157 3796 5648 3846
rect 4099 3778 4157 3788
rect 5706 3796 6163 3846
rect 5648 3778 5706 3788
rect 6163 3778 6221 3788
rect 6287 3819 6384 3937
rect 6287 3741 6297 3819
rect 6377 3741 6384 3819
rect 6287 3731 6384 3741
rect -7751 -848 -7631 3708
rect -3159 3668 -3033 3708
rect 2551 3678 5189 3688
rect -4931 3658 -1261 3668
rect -4873 3600 -1319 3658
rect 2609 3628 3067 3678
rect 2551 3610 2609 3620
rect 3125 3628 4615 3678
rect 3067 3610 3125 3620
rect 4673 3628 5131 3678
rect 4615 3610 4673 3620
rect 5131 3610 5189 3620
rect -4931 3590 -1261 3600
rect 2809 2435 2867 2445
rect 4873 2435 4931 2445
rect 2867 2377 4873 2397
rect 4931 2377 7354 2397
rect 2809 2337 7354 2377
rect 7114 2239 7194 2257
rect -6109 2165 -6017 2184
rect -6109 2107 -6094 2165
rect -6036 2107 -6017 2165
rect 7114 2181 7125 2239
rect 7183 2181 7194 2239
rect -6109 2097 6625 2107
rect -6612 2064 -6554 2065
rect -6625 2055 -6533 2064
rect -6625 1997 -6612 2055
rect -6554 1997 -6533 2055
rect -6017 2037 -5851 2097
rect -5759 2037 -5077 2097
rect -4985 2037 -4819 2097
rect -4727 2037 -4045 2097
rect -3953 2037 -3787 2097
rect -3695 2037 -3013 2097
rect -2921 2037 -2755 2097
rect -2663 2037 -1981 2097
rect -1889 2037 -1723 2097
rect -1631 2037 -949 2097
rect -857 2037 -691 2097
rect -599 2037 341 2097
rect 433 2037 1115 2097
rect 1207 2037 1373 2097
rect 1465 2037 2147 2097
rect 2239 2037 2405 2097
rect 2497 2037 3179 2097
rect 3271 2037 3437 2097
rect 3529 2037 4211 2097
rect 4303 2037 4469 2097
rect 4561 2037 5243 2097
rect 5335 2037 5501 2097
rect 5593 2037 6275 2097
rect 6367 2037 6533 2097
rect -6109 2027 6625 2037
rect -6625 1987 -6533 1997
rect -6625 1977 6109 1987
rect -6533 1917 -6367 1977
rect -6275 1917 -5593 1977
rect -5501 1917 -5335 1977
rect -5243 1917 -4561 1977
rect -4469 1917 -4303 1977
rect -4211 1917 -3529 1977
rect -3437 1917 -3271 1977
rect -3179 1917 -2497 1977
rect -2405 1917 -2239 1977
rect -2147 1917 -1465 1977
rect -1373 1917 -1207 1977
rect -1115 1917 -433 1977
rect -341 1917 599 1977
rect 691 1917 857 1977
rect 949 1917 1631 1977
rect 1723 1917 1889 1977
rect 1981 1917 2663 1977
rect 2755 1917 2921 1977
rect 3013 1917 3695 1977
rect 3787 1917 3953 1977
rect 4045 1917 4727 1977
rect 4819 1917 4985 1977
rect 5077 1917 5759 1977
rect 5851 1917 6017 1977
rect -6625 1907 6109 1917
rect -5963 700 6479 710
rect -5905 642 -4931 700
rect -4873 642 -3899 700
rect -3841 642 -2867 700
rect -2809 642 -1835 700
rect -1777 642 -803 700
rect -745 642 229 700
rect 287 642 1261 700
rect 1319 642 2293 700
rect 2351 642 3325 700
rect 3383 642 4357 700
rect 4415 642 5389 700
rect 5447 642 6421 700
rect -5963 632 6479 642
rect -3383 570 -3325 571
rect 745 570 803 571
rect -6479 561 5963 570
rect -6479 560 -3383 561
rect -6421 502 -5447 560
rect -5389 502 -4415 560
rect -4357 503 -3383 560
rect -3325 560 745 561
rect -3325 503 -2351 560
rect -4357 502 -2351 503
rect -2293 502 -1319 560
rect -1261 502 -287 560
rect -229 503 745 560
rect 803 560 5963 561
rect 803 503 1777 560
rect -229 502 1777 503
rect 1835 502 2809 560
rect 2867 502 3841 560
rect 3899 502 4873 560
rect 4931 502 5905 560
rect -6479 492 5963 502
rect -298 -320 -218 492
rect -298 -378 -287 -320
rect -229 -378 -218 -320
rect -298 -388 -218 -378
rect -29 401 29 411
rect -29 -320 29 343
rect -29 -392 29 -378
rect 218 401 298 411
rect 218 343 229 401
rect 287 343 298 401
rect 218 -320 298 343
rect 218 -378 229 -320
rect 287 -378 298 -320
rect 218 -389 298 -378
rect 7114 -458 7194 2181
rect 7274 -59 7354 2337
rect -555 -538 7194 -458
rect 7275 -433 7354 -59
rect 7275 -443 7475 -433
rect -555 -578 -477 -538
rect 7275 -578 7377 -443
rect -1577 -588 545 -578
rect -1519 -646 487 -588
rect -1577 -656 545 -646
rect 616 -588 7377 -578
rect 674 -643 7377 -588
rect 674 -646 7475 -643
rect 616 -656 7475 -646
rect -3899 -706 3383 -696
rect -3841 -764 -2867 -706
rect -2809 -764 -1835 -706
rect -1777 -764 -1319 -706
rect -1261 -764 229 -706
rect 287 -764 745 -706
rect 803 -764 2293 -706
rect 2351 -764 3325 -706
rect -3899 -774 3383 -764
rect -545 -824 1577 -814
rect -7751 -968 -5708 -848
rect -487 -825 1519 -824
rect -487 -882 616 -825
rect -545 -883 616 -882
rect 674 -882 1519 -825
rect 674 -883 1577 -882
rect -545 -892 1577 -883
rect 616 -893 674 -892
rect -5828 -2390 -5708 -968
rect -3383 -942 3899 -932
rect -3325 -1000 -2351 -942
rect -2293 -1000 -803 -942
rect -745 -1000 -287 -942
rect -229 -1000 1261 -942
rect 1319 -1000 1777 -942
rect 1835 -1000 2809 -942
rect 2867 -1000 3841 -942
rect -3383 -1010 3899 -1000
rect -4415 -2130 -4357 -2120
rect -4415 -2228 -4357 -2188
rect 4357 -2130 4415 -2120
rect 4357 -2228 4415 -2188
rect -4415 -2328 4415 -2228
rect -50 -2390 50 -2328
rect -5828 -2490 50 -2390
rect 255 -2444 313 -2434
rect 255 -2512 313 -2502
rect -8756 -3956 -8156 -3946
rect -8756 -4266 -8156 -4256
rect 8156 -3956 8756 -3946
rect 8156 -4266 8756 -4256
<< via2 >>
rect -8756 3956 -8156 4256
rect 8156 3956 8756 4256
rect -2349 3784 -2291 3842
rect 6297 3741 6377 3819
rect -6094 2107 -6036 2165
rect -6612 1997 -6554 2055
rect 7377 -643 7475 -443
rect 255 -2502 313 -2444
rect -8756 -4256 -8156 -3956
rect 8156 -4256 8756 -3956
<< metal3 >>
rect -8766 4256 -8146 4261
rect -8766 3956 -8756 4256
rect -8156 3956 -8146 4256
rect 8146 4256 8766 4261
rect -8766 3951 -8146 3956
rect 3150 3934 7096 4034
rect 8146 3956 8156 4256
rect 8756 3956 8766 4256
rect 8146 3951 8766 3956
rect 3150 3867 3250 3934
rect -2362 3842 3250 3867
rect -2362 3784 -2349 3842
rect -2291 3784 3250 3842
rect -2362 3767 3250 3784
rect 6287 3819 6902 3826
rect 6287 3741 6297 3819
rect 6377 3741 6902 3819
rect 6287 3731 6902 3741
rect 6807 2562 6902 3731
rect 6996 2933 7096 3934
rect 6996 2833 8433 2933
rect 6807 2467 8064 2562
rect -7967 2250 -6259 2350
rect -7967 141 -7867 2250
rect -6359 2202 -6259 2250
rect -6359 2165 -6026 2202
rect -6359 2107 -6094 2165
rect -6036 2107 -6026 2165
rect -6359 2102 -6026 2107
rect 7969 2187 8064 2467
rect 8333 2418 8433 2833
rect 8333 2403 9359 2418
rect 8334 2318 9359 2403
rect -8536 41 -7867 141
rect -7404 2055 -6544 2092
rect 7969 2087 9359 2187
rect -7404 1997 -6612 2055
rect -6554 1997 -6544 2055
rect -7404 1992 -6544 1997
rect -7404 -104 -7304 1992
rect -8545 -204 -7304 -104
rect 7745 -110 14758 90
rect 7367 -443 7485 -438
rect 7745 -443 7945 -110
rect 7367 -643 7377 -443
rect 7475 -643 7945 -443
rect 8339 -580 9359 -480
rect 7367 -648 7485 -643
rect 8339 -2426 8439 -580
rect 233 -2444 8439 -2426
rect 233 -2502 255 -2444
rect 313 -2502 8439 -2444
rect 233 -2526 8439 -2502
rect -8542 -2942 9499 -2742
rect -8766 -3956 -8146 -3951
rect -8766 -4256 -8756 -3956
rect -8156 -4256 -8146 -3956
rect -8766 -4261 -8146 -4256
rect 8146 -3956 8766 -3951
rect 8146 -4256 8156 -3956
rect 8756 -4256 8766 -3956
rect 8146 -4261 8766 -4256
<< via3 >>
rect -8756 3956 -8156 4256
rect 8156 3956 8756 4256
rect -8756 -4256 -8156 -3956
rect 8156 -4256 8756 -3956
<< metal4 >>
rect -9000 4256 9000 4500
rect -9000 3956 -8756 4256
rect -8156 3956 8156 4256
rect 8756 3956 9000 4256
rect -9000 3700 9000 3956
rect -9000 -3956 9000 -3700
rect -9000 -4256 -8756 -3956
rect -8156 -4256 8156 -3956
rect 8756 -4256 9000 -3956
rect -9000 -4500 9000 -4256
<< comment >>
rect -3111 2071 -3087 2248
rect 4375 1995 4394 2140
rect -19 -187 18 122
use cascode_bias  cascode_bias_0
timestamp 1624430562
transform 1 0 12000 0 1 0
box -3000 -4500 3000 4500
use sky130_fd_pr__pfet_g5v0d10v5_QM5ZLW  xm4
timestamp 1624430562
transform 1 0 4386 0 1 3000
box -2417 -600 2417 600
use sky130_fd_pr__pfet_g5v0d10v5_QF5B2D  xm2
timestamp 1624430562
transform 1 0 0 0 1 1300
box -7061 -600 7061 600
use sky130_fd_pr__nfet_g5v0d10v5_V3Y342  xm1
timestamp 1624430562
transform 1 0 0 0 1 -1600
box -4673 -588 4673 588
use sky130_fd_pr__pfet_g5v0d10v5_QC2ZLW  xm3
timestamp 1624430562
transform 1 0 -3096 0 1 3000
box -2159 -600 2159 600
<< labels >>
flabel metal4 -9000 3700 -9000 4500 3 FreeSans 480 0 0 0 vdd
port 5 e
flabel metal4 -9000 -4500 -9000 -3700 3 FreeSans 480 0 0 0 vss
port 6 e
flabel metal3 14758 -110 14758 90 1 FreeSans 240 0 0 0 out
port 4 n
flabel metal3 -8542 -2941 -8541 -2742 1 FreeSans 240 0 0 0 ibias
port 1 n
flabel metal3 -8536 41 -8536 141 1 FreeSans 240 0 0 0 in_p
port 3 n
flabel metal3 -8545 -204 -8544 -104 1 FreeSans 240 0 0 0 in_m
port 2 n
<< properties >>
string FIXED_BBOX -8842 -4342 8842 -198
<< end >>
