magic
tech sky130A
magscale 1 2
timestamp 1384693831
<< checkpaint >>
rect -1378 -1378 3746 3948
<< metal1 >>
rect 570 1034 1838 1036
rect 570 982 576 1034
rect 628 982 1780 1034
rect 1832 982 1838 1034
rect 570 980 1838 982
rect 656 278 1752 280
rect 656 226 662 278
rect 714 226 1694 278
rect 1746 226 1752 278
rect 656 224 1752 226
<< via1 >>
rect 576 982 628 1034
rect 1780 982 1832 1034
rect 662 226 714 278
rect 1694 226 1746 278
<< metal2 >>
rect 1864 1792 1920 1801
rect 1864 1727 1920 1736
rect 574 1034 630 1040
rect 574 982 576 1034
rect 628 982 630 1034
rect 574 976 630 982
rect 1778 1034 1834 1040
rect 1778 982 1780 1034
rect 1832 982 1834 1034
rect 1778 976 1834 982
rect 488 280 544 289
rect 488 215 544 224
rect 660 278 716 284
rect 660 226 662 278
rect 714 226 716 278
rect 660 220 716 226
rect 1692 278 1748 284
rect 1692 226 1694 278
rect 1746 226 1748 278
rect 1692 220 1748 226
<< via2 >>
rect 1864 1736 1920 1792
rect 488 224 544 280
<< metal3 >>
rect -80 1796 2448 1844
rect -80 1792 2336 1796
rect -80 1736 1864 1792
rect 1920 1736 2336 1792
rect -80 1732 2336 1736
rect 2400 1732 2448 1796
rect -80 1684 2448 1732
rect 483 284 625 332
rect 483 280 560 284
rect 483 224 488 280
rect 544 224 560 280
rect 483 220 560 224
rect 624 220 625 284
rect 483 172 625 220
rect -80 32 2448 80
rect -80 -32 -32 32
rect 32 -32 560 32
rect 624 -32 2448 32
rect -80 -80 2448 -32
<< via3 >>
rect 2336 1732 2400 1796
rect 560 220 624 284
rect -32 -32 32 32
rect 560 -32 624 32
<< metal4 >>
rect -118 32 118 1882
rect 2250 1796 2486 1882
rect 2250 1732 2336 1796
rect 2400 1732 2486 1796
rect -118 -32 -32 32
rect 32 -32 118 32
rect -118 -118 118 -32
rect 474 284 710 285
rect 474 220 560 284
rect 624 220 710 284
rect 474 32 710 220
rect 474 -32 560 32
rect 624 -32 710 32
rect 474 -33 710 -32
rect 2250 -118 2486 1732
use NMOS_S_6078655_X5_Y2_1678793193  NMOS_S_6078655_X5_Y2_1678793193_0
timestamp 1374899056
transform 1 0 1204 0 1 0
box 121 52 1083 2658
use PMOS_S_79543009_X5_Y2_1678793194  PMOS_S_79543009_X5_Y2_1678793194_0
timestamp 1374899056
transform -1 0 1204 0 1 0
box 0 0 1204 2688
<< labels >>
flabel metal2 s 688 672 688 672 0 FreeSerif 0 0 0 0 Y
flabel metal2 s 602 1512 602 1512 0 FreeSerif 0 0 0 0 A
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal3 s 554 252 554 252 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
<< end >>
