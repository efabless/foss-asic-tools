magic
tech sky130A
magscale 1 2
timestamp 1620965225
<< error_p >>
rect -29 581 29 587
rect -29 547 -17 581
rect -29 541 29 547
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect -29 -587 29 -581
<< nwell >>
rect -308 -797 308 797
<< mvpmos >>
rect -50 -500 50 500
<< mvpdiff >>
rect -108 488 -50 500
rect -108 -488 -96 488
rect -62 -488 -50 488
rect -108 -500 -50 -488
rect 50 488 108 500
rect 50 -488 62 488
rect 96 -488 108 488
rect 50 -500 108 -488
<< mvpdiffc >>
rect -96 -488 -62 488
rect 62 -488 96 488
<< mvnsubdiff >>
rect -242 719 242 731
rect -242 685 -134 719
rect 134 685 242 719
rect -242 673 242 685
rect -242 623 -184 673
rect -242 -623 -230 623
rect -196 -623 -184 623
rect 184 623 242 673
rect -242 -673 -184 -623
rect 184 -623 196 623
rect 230 -623 242 623
rect 184 -673 242 -623
rect -242 -685 242 -673
rect -242 -719 -134 -685
rect 134 -719 242 -685
rect -242 -731 242 -719
<< mvnsubdiffcont >>
rect -134 685 134 719
rect -230 -623 -196 623
rect 196 -623 230 623
rect -134 -719 134 -685
<< poly >>
rect -50 581 50 597
rect -50 547 -34 581
rect 34 547 50 581
rect -50 500 50 547
rect -50 -547 50 -500
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -597 50 -581
<< polycont >>
rect -34 547 34 581
rect -34 -581 34 -547
<< locali >>
rect -230 685 -134 719
rect 134 685 230 719
rect -230 623 -196 685
rect 196 623 230 685
rect -50 547 -34 581
rect 34 547 50 581
rect -96 488 -62 504
rect -96 -504 -62 -488
rect 62 488 96 504
rect 62 -504 96 -488
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -230 -685 -196 -623
rect 196 -685 230 -623
rect -230 -719 -134 -685
rect 134 -719 230 -685
<< viali >>
rect -17 547 17 581
rect -96 -488 -62 488
rect 62 -488 96 488
rect -17 -581 17 -547
<< metal1 >>
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect -102 488 -56 500
rect -102 -488 -96 488
rect -62 -488 -56 488
rect -102 -500 -56 -488
rect 56 488 102 500
rect 56 -488 62 488
rect 96 -488 102 488
rect 56 -500 102 -488
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -213 -702 213 702
string parameters w 5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
