magic
tech sky130A
magscale 1 2
timestamp 1622253817
<< nwell >>
rect -11400 5300 6900 9000
rect -11400 1000 -4600 5300
rect -11723 -4877 -11623 -4763
<< pwell >>
rect -4500 0 6900 5100
<< mvpsubdiff >>
rect -4434 5022 6834 5034
rect -4434 4862 -4200 5022
rect 6600 4862 6834 5022
rect -4434 4850 6834 4862
rect -4434 4800 -4250 4850
rect -4434 300 -4422 4800
rect -4262 300 -4250 4800
rect -4434 250 -4250 300
rect 6650 4800 6834 4850
rect 6650 300 6662 4800
rect 6822 300 6834 4800
rect 6650 250 6834 300
rect -4434 238 6834 250
rect -4434 78 -4200 238
rect 6600 78 6834 238
rect -4434 66 6834 78
<< mvnsubdiff >>
rect -11334 8922 -4666 8934
rect -11334 8762 -11100 8922
rect -4900 8762 -4666 8922
rect -11334 8750 -4666 8762
rect -11334 8700 -11150 8750
rect -11334 1300 -11322 8700
rect -11162 1300 -11150 8700
rect -11334 1250 -11150 1300
rect -4850 8700 -4666 8750
rect -4850 1300 -4838 8700
rect -4678 1300 -4666 8700
rect -4434 8922 6834 8934
rect -4434 8762 -4200 8922
rect 6600 8762 6834 8922
rect -4434 8750 6834 8762
rect -4434 8700 -4250 8750
rect -4434 5600 -4422 8700
rect -4262 5600 -4250 8700
rect -4434 5550 -4250 5600
rect 6650 8700 6834 8750
rect 6650 5600 6662 8700
rect 6822 5600 6834 8700
rect 6650 5550 6834 5600
rect -4434 5538 6834 5550
rect -4434 5378 -4200 5538
rect 6600 5378 6834 5538
rect -4434 5366 6834 5378
rect -4850 1250 -4666 1300
rect -11334 1238 -4666 1250
rect -11334 1078 -11100 1238
rect -4900 1078 -4666 1238
rect -11334 1066 -4666 1078
<< mvpsubdiffcont >>
rect -4200 4862 6600 5022
rect -4422 300 -4262 4800
rect 6662 300 6822 4800
rect -4200 78 6600 238
<< mvnsubdiffcont >>
rect -11100 8762 -4900 8922
rect -11322 1300 -11162 8700
rect -4838 1300 -4678 8700
rect -4200 8762 6600 8922
rect -4422 5600 -4262 8700
rect 6662 5600 6822 8700
rect -4200 5378 6600 5538
rect -11100 1078 -4900 1238
<< locali >>
rect -11322 8700 -11162 8922
rect -11322 1078 -11162 1300
rect -4838 8700 -4678 8922
rect -4422 8700 -4262 8922
rect -4422 5378 -4262 5600
rect 6662 8700 6822 8922
rect 6662 5378 6822 5600
rect -4838 1078 -4678 1300
rect -4422 4800 -4262 5022
rect -4422 78 -4262 300
rect 6662 4800 6822 5022
rect 6662 78 6822 300
<< viali >>
rect -11162 8762 -11100 8922
rect -11100 8762 -4900 8922
rect -4900 8762 -4838 8922
rect -11322 1614 -11162 8386
rect -4838 1614 -4678 8386
rect -4262 8762 -4200 8922
rect -4200 8762 6600 8922
rect 6600 8762 6662 8922
rect -4422 5699 -4262 8601
rect 6662 5699 6822 8601
rect -4262 5378 -4200 5538
rect -4200 5378 6600 5538
rect 6600 5378 6662 5538
rect -11162 1078 -11100 1238
rect -11100 1078 -4900 1238
rect -4900 1078 -4838 1238
rect -4262 4862 -4200 5022
rect -4200 4862 6600 5022
rect 6600 4862 6662 5022
rect -4422 469 -4262 4631
rect 6662 469 6822 4631
rect -4262 78 -4200 238
rect -4200 78 6600 238
rect 6600 78 6662 238
<< metal1 >>
rect -11328 8922 -4672 8928
rect -11328 8762 -11162 8922
rect -4838 8762 -4672 8922
rect -11328 8756 -4672 8762
rect -11328 8386 -11156 8756
rect -10556 8456 -10546 8756
rect -5454 8456 -5444 8756
rect -11328 1614 -11322 8386
rect -11162 1614 -11156 8386
rect -11328 1244 -11156 1614
rect -4844 8386 -4672 8756
rect -4844 1614 -4838 8386
rect -4678 1614 -4672 8386
rect -4428 8922 6828 8928
rect -4428 8762 -4262 8922
rect 6662 8762 6828 8922
rect -4428 8756 6828 8762
rect -4428 8601 -4256 8756
rect -4428 5699 -4422 8601
rect -4262 8456 -4256 8601
rect -3656 8456 6056 8756
rect 6656 8601 6828 8756
rect 6656 8456 6662 8601
rect -4262 8200 6662 8456
rect -4262 5699 -4256 8200
rect 2571 7690 2921 8200
rect 4225 7690 4575 8200
rect 5879 7690 6229 8200
rect -3661 7671 2061 7690
rect -3661 7468 -3641 7671
rect -3417 7468 2061 7671
rect -3661 7450 2061 7468
rect -3661 7337 -3615 7450
rect -3403 7337 -3357 7450
rect -3145 7337 -3099 7450
rect -2887 7337 -2841 7450
rect -2629 7337 -2583 7450
rect -2371 7337 -2325 7450
rect -3661 7291 -2325 7337
rect -3661 7250 -3615 7291
rect -3403 7250 -3357 7291
rect -3145 7250 -3099 7291
rect -2887 7250 -2841 7291
rect -2629 7250 -2583 7291
rect -2371 7250 -2325 7291
rect -1855 7250 -1809 7450
rect -1339 7250 -1293 7450
rect -823 7250 -777 7450
rect -307 7250 -261 7450
rect 209 7250 255 7450
rect 725 7337 771 7450
rect 983 7337 1029 7450
rect 1241 7337 1287 7450
rect 1499 7337 1545 7450
rect 1757 7337 1803 7450
rect 2015 7337 2061 7450
rect 725 7291 2061 7337
rect 725 7250 771 7291
rect 983 7250 1029 7291
rect 1241 7250 1287 7291
rect 1499 7250 1545 7291
rect 1757 7250 1803 7291
rect 2015 7250 2061 7291
rect 2571 7450 6229 7690
rect 2571 7337 2617 7450
rect 2829 7337 2875 7450
rect 2571 7291 2875 7337
rect 2571 7250 2617 7291
rect 2829 7250 2875 7291
rect 3345 7250 3391 7450
rect 3861 7250 3907 7450
rect 4377 7250 4423 7450
rect 4893 7250 4939 7450
rect 5409 7250 5455 7450
rect 5925 7337 5971 7450
rect 6183 7337 6229 7450
rect 5925 7291 6229 7337
rect 5925 7250 5971 7291
rect 6183 7250 6229 7291
rect -2265 6149 -2173 6163
rect -2265 6123 -2245 6149
rect -2255 6097 -2245 6123
rect -2193 6123 -2173 6149
rect -2193 6097 -2183 6123
rect -2113 6050 -2067 6250
rect -2007 6149 -1915 6163
rect -2007 6123 -1987 6149
rect -1997 6097 -1987 6123
rect -1935 6123 -1915 6149
rect -1749 6149 -1657 6163
rect -1749 6123 -1729 6149
rect -1935 6097 -1925 6123
rect -1739 6097 -1729 6123
rect -1677 6123 -1657 6149
rect -1677 6097 -1667 6123
rect -1597 6050 -1551 6250
rect -1491 6149 -1399 6163
rect -1491 6123 -1471 6149
rect -1481 6097 -1471 6123
rect -1419 6123 -1399 6149
rect -1233 6149 -1141 6163
rect -1233 6123 -1213 6149
rect -1419 6097 -1409 6123
rect -1223 6097 -1213 6123
rect -1161 6123 -1141 6149
rect -1161 6097 -1151 6123
rect -1081 6050 -1035 6250
rect -975 6149 -883 6163
rect -975 6123 -955 6149
rect -965 6097 -955 6123
rect -903 6123 -883 6149
rect -717 6149 -625 6163
rect -717 6123 -697 6149
rect -903 6097 -893 6123
rect -707 6097 -697 6123
rect -645 6123 -625 6149
rect -645 6097 -635 6123
rect -565 6050 -519 6250
rect -459 6149 -367 6163
rect -459 6123 -439 6149
rect -449 6097 -439 6123
rect -387 6123 -367 6149
rect -201 6149 -109 6163
rect -201 6123 -181 6149
rect -387 6097 -377 6123
rect -191 6097 -181 6123
rect -129 6123 -109 6149
rect -129 6097 -119 6123
rect -49 6050 -3 6250
rect 57 6149 149 6163
rect 57 6123 77 6149
rect 67 6097 77 6123
rect 129 6123 149 6149
rect 315 6149 407 6163
rect 315 6123 335 6149
rect 129 6097 139 6123
rect 325 6097 335 6123
rect 387 6123 407 6149
rect 387 6097 397 6123
rect 467 6050 513 6250
rect 3087 6209 3133 6250
rect 2935 6163 3543 6209
rect 573 6149 665 6163
rect 573 6123 593 6149
rect 583 6097 593 6123
rect 645 6123 665 6149
rect 645 6097 655 6123
rect -2113 6035 513 6050
rect -2113 5835 -900 6035
rect -700 5835 513 6035
rect -2113 5810 513 5835
rect 3050 5893 3170 6163
rect 3603 6036 3649 6250
rect 4119 6209 4165 6250
rect 4635 6209 4681 6250
rect 3709 6163 5091 6209
rect 3590 5984 3600 6036
rect 3652 5984 3662 6036
rect 4082 5893 4202 6163
rect 4598 5893 4718 6163
rect 5151 6036 5197 6250
rect 5667 6209 5713 6250
rect 5257 6163 5865 6209
rect 5138 5984 5148 6036
rect 5200 5984 5210 6036
rect 5630 5893 5750 6163
rect 3050 5813 5750 5893
rect 3050 5733 4320 5813
rect -4428 5544 -4256 5699
rect 4310 5653 4320 5733
rect 4480 5733 5750 5813
rect 4480 5653 4490 5733
rect 6656 5699 6662 8200
rect 6822 5699 6828 8601
rect 7835 7848 9946 7926
rect 7835 7802 9627 7848
rect 7835 7642 7868 7802
rect 8028 7642 9627 7802
rect 7835 7605 9627 7642
rect 9867 7605 9946 7848
rect 7835 7506 9946 7605
rect 7835 7505 9531 7506
rect 6656 5544 6828 5699
rect -4428 5538 6828 5544
rect -4428 5378 -4262 5538
rect 6662 5378 6828 5538
rect -4428 5372 6828 5378
rect -4844 1244 -4672 1614
rect -11328 1238 -4672 1244
rect -11328 1078 -11162 1238
rect -4838 1078 -4672 1238
rect -11328 1072 -4672 1078
rect -4428 5022 6828 5028
rect -4428 4862 -4262 5022
rect 6662 4862 6828 5022
rect -4428 4856 6828 4862
rect -4428 4631 -4256 4856
rect -4428 469 -4422 4631
rect -4262 800 -4256 4631
rect -1745 4625 2945 4640
rect -1745 4425 500 4625
rect 700 4425 2945 4625
rect -1745 4400 2945 4425
rect -1745 4178 -1699 4400
rect -1242 4314 -1232 4366
rect -1180 4314 -1170 4366
rect -1897 4132 -1289 4178
rect -1745 4100 -1699 4132
rect -1229 4100 -1183 4314
rect -713 4178 -667 4400
rect -210 4314 -200 4366
rect -148 4314 -138 4366
rect -1123 4132 -257 4178
rect -713 4100 -667 4132
rect -197 4100 -151 4314
rect 319 4178 365 4400
rect 835 4178 881 4400
rect 1338 4314 1348 4366
rect 1400 4314 1410 4366
rect -91 4132 1291 4178
rect 319 4100 365 4132
rect 835 4100 881 4132
rect 1351 4100 1397 4314
rect 1867 4178 1913 4400
rect 2370 4314 2380 4366
rect 2432 4314 2442 4366
rect 1457 4132 2323 4178
rect 1867 4100 1913 4132
rect 2383 4100 2429 4314
rect 2899 4178 2945 4400
rect 6656 4631 6828 4856
rect 2489 4132 3097 4178
rect 2899 4100 2945 4132
rect -3293 3068 -3247 3100
rect -3035 3068 -2989 3100
rect -2777 3068 -2731 3100
rect -2519 3068 -2473 3100
rect -2261 3068 -2215 3100
rect -2003 3068 -1957 3100
rect -1745 3068 -1699 3100
rect -3293 3022 -1957 3068
rect -1897 3048 -1547 3068
rect -1897 3022 -1748 3048
rect -3293 2900 -3247 3022
rect -3035 2900 -2989 3022
rect -2777 2900 -2731 3022
rect -2519 2900 -2473 3022
rect -2261 2900 -2215 3022
rect -2003 2900 -1957 3022
rect -1758 2996 -1748 3022
rect -1696 3022 -1547 3048
rect -1696 2996 -1686 3022
rect -1487 2900 -1441 3100
rect -971 2900 -925 3100
rect -713 3068 -667 3100
rect -865 3048 -515 3068
rect -865 3022 -716 3048
rect -726 2996 -716 3022
rect -664 3022 -515 3048
rect -664 2996 -654 3022
rect -455 2900 -409 3100
rect 61 2900 107 3100
rect 319 3068 365 3100
rect 167 3048 517 3068
rect 167 3022 316 3048
rect 306 2996 316 3022
rect 368 3022 517 3048
rect 368 2996 378 3022
rect 577 2900 623 3100
rect 835 3068 881 3100
rect 683 3048 1033 3068
rect 683 3022 832 3048
rect 822 2996 832 3022
rect 884 3022 1033 3048
rect 884 2996 894 3022
rect 1093 2900 1139 3100
rect 1609 2900 1655 3100
rect 1867 3068 1913 3100
rect 1715 3048 2065 3068
rect 1715 3022 1864 3048
rect 1854 2996 1864 3022
rect 1916 3022 2065 3048
rect 1916 2996 1926 3022
rect 2125 2900 2171 3100
rect 2641 2900 2687 3100
rect 2899 3068 2945 3100
rect 3157 3068 3203 3100
rect 3415 3068 3461 3100
rect 3673 3068 3719 3100
rect 3931 3068 3977 3100
rect 4189 3068 4235 3100
rect 4447 3068 4493 3100
rect 2747 3048 3097 3068
rect 2747 3022 2896 3048
rect 2886 2996 2896 3022
rect 2948 3022 3097 3048
rect 3157 3022 4493 3068
rect 2948 2996 2958 3022
rect 3157 2900 3203 3022
rect 3415 2900 3461 3022
rect 3673 2900 3719 3022
rect 3931 2900 3977 3022
rect 4189 2900 4235 3022
rect 4447 2900 4493 3022
rect -3293 2500 4493 2900
rect -3293 800 -2361 2500
rect -1745 2450 3398 2460
rect -1745 2210 3148 2450
rect 3388 2210 3398 2450
rect -1745 2200 3398 2210
rect -1887 2112 -1877 2138
rect -1897 2086 -1877 2112
rect -1825 2112 -1815 2138
rect -1825 2086 -1805 2112
rect -1897 2078 -1805 2086
rect -1745 2000 -1699 2200
rect -1629 2112 -1619 2138
rect -1639 2086 -1619 2112
rect -1567 2112 -1557 2138
rect -1371 2112 -1361 2138
rect -1567 2086 -1547 2112
rect -1639 2078 -1547 2086
rect -1381 2086 -1361 2112
rect -1309 2112 -1299 2138
rect -1309 2086 -1289 2112
rect -1381 2078 -1289 2086
rect -1229 2000 -1183 2200
rect -1113 2112 -1103 2138
rect -1123 2086 -1103 2112
rect -1051 2112 -1041 2138
rect -855 2112 -845 2138
rect -1051 2086 -1031 2112
rect -1123 2078 -1031 2086
rect -865 2086 -845 2112
rect -793 2112 -783 2138
rect -793 2086 -773 2112
rect -865 2078 -773 2086
rect -713 2000 -667 2200
rect -597 2112 -587 2138
rect -607 2086 -587 2112
rect -535 2112 -525 2138
rect -339 2112 -329 2138
rect -535 2086 -515 2112
rect -607 2078 -515 2086
rect -349 2086 -329 2112
rect -277 2112 -267 2138
rect -277 2086 -257 2112
rect -349 2078 -257 2086
rect -197 2000 -151 2200
rect -81 2112 -71 2138
rect -91 2086 -71 2112
rect -19 2112 -9 2138
rect 177 2112 187 2138
rect -19 2086 1 2112
rect -91 2078 1 2086
rect 167 2086 187 2112
rect 239 2112 249 2138
rect 239 2086 259 2112
rect 167 2078 259 2086
rect 319 2000 365 2200
rect 435 2112 445 2138
rect 425 2086 445 2112
rect 497 2112 507 2138
rect 693 2112 703 2138
rect 497 2086 517 2112
rect 425 2032 517 2086
rect 683 2086 703 2112
rect 755 2112 765 2138
rect 755 2086 775 2112
rect 683 2078 775 2086
rect 835 2000 881 2200
rect 951 2112 961 2138
rect 941 2086 961 2112
rect 1013 2112 1023 2138
rect 1209 2112 1219 2138
rect 1013 2086 1033 2112
rect 941 2078 1033 2086
rect 1199 2086 1219 2112
rect 1271 2112 1281 2138
rect 1271 2086 1291 2112
rect 1199 2078 1291 2086
rect 1351 2000 1397 2200
rect 1467 2112 1477 2138
rect 1457 2086 1477 2112
rect 1529 2112 1539 2138
rect 1725 2112 1735 2138
rect 1529 2086 1549 2112
rect 1457 2078 1549 2086
rect 1715 2086 1735 2112
rect 1787 2112 1797 2138
rect 1787 2086 1807 2112
rect 1715 2078 1807 2086
rect 1867 2000 1913 2200
rect 1983 2112 1993 2138
rect 1973 2086 1993 2112
rect 2045 2112 2055 2138
rect 2241 2112 2251 2138
rect 2045 2086 2065 2112
rect 1973 2078 2065 2086
rect 2231 2086 2251 2112
rect 2303 2112 2313 2138
rect 2303 2086 2323 2112
rect 2231 2078 2323 2086
rect 2383 2000 2429 2200
rect 2499 2112 2509 2138
rect 2489 2086 2509 2112
rect 2561 2112 2571 2138
rect 2757 2112 2767 2138
rect 2561 2086 2581 2112
rect 2489 2078 2581 2086
rect 2747 2086 2767 2112
rect 2819 2112 2829 2138
rect 2819 2086 2839 2112
rect 2747 2078 2839 2086
rect 2899 2000 2945 2200
rect 3015 2112 3025 2138
rect 3005 2086 3025 2112
rect 3077 2112 3087 2138
rect 3077 2086 3097 2112
rect 3005 2078 3097 2086
rect -2261 968 -2215 1000
rect -2003 968 -1957 1000
rect -2261 922 -1957 968
rect -2261 800 -2215 922
rect -2003 800 -1957 922
rect -1487 800 -1441 1000
rect -971 800 -925 1000
rect -455 800 -409 1000
rect 61 800 107 1000
rect 577 800 623 1000
rect 1093 800 1139 1000
rect 1609 800 1655 1000
rect 2125 800 2171 1000
rect 2641 800 2687 1000
rect 3157 968 3203 1000
rect 3415 968 3461 1000
rect 3157 922 3461 968
rect 3157 800 3203 922
rect 3415 800 3461 922
rect 3561 800 4493 2500
rect 6656 800 6662 4631
rect -4262 544 6662 800
rect -4262 469 -4256 544
rect -4428 244 -4256 469
rect -3656 244 6056 544
rect 6656 469 6662 544
rect 6822 469 6828 4631
rect 6656 244 6828 469
rect -4428 238 6828 244
rect -4428 78 -4262 238
rect 6662 78 6828 238
rect -4428 72 6828 78
rect 8066 634 9531 1495
rect 8066 85 8369 634
rect 9186 85 9531 634
rect 8066 4 9531 85
<< via1 >>
rect -11156 8456 -10556 8756
rect -5444 8456 -4844 8756
rect -4256 8456 -3656 8756
rect 6056 8456 6656 8756
rect -3641 7468 -3417 7671
rect -2245 6097 -2193 6149
rect -1987 6097 -1935 6149
rect -1729 6097 -1677 6149
rect -1471 6097 -1419 6149
rect -1213 6097 -1161 6149
rect -955 6097 -903 6149
rect -697 6097 -645 6149
rect -439 6097 -387 6149
rect -181 6097 -129 6149
rect 77 6097 129 6149
rect 335 6097 387 6149
rect 593 6097 645 6149
rect -900 5835 -700 6035
rect 3600 5984 3652 6036
rect 5148 5984 5200 6036
rect 4320 5653 4480 5813
rect 7868 7642 8028 7802
rect 9627 7605 9867 7848
rect 500 4425 700 4625
rect -1232 4314 -1180 4366
rect -200 4314 -148 4366
rect 1348 4314 1400 4366
rect 2380 4314 2432 4366
rect -1748 2996 -1696 3048
rect -716 2996 -664 3048
rect 316 2996 368 3048
rect 832 2996 884 3048
rect 1864 2996 1916 3048
rect 2896 2996 2948 3048
rect 3148 2210 3388 2450
rect -1877 2086 -1825 2138
rect -1619 2086 -1567 2138
rect -1361 2086 -1309 2138
rect -1103 2086 -1051 2138
rect -845 2086 -793 2138
rect -587 2086 -535 2138
rect -329 2086 -277 2138
rect -71 2086 -19 2138
rect 187 2086 239 2138
rect 445 2086 497 2138
rect 703 2086 755 2138
rect 961 2086 1013 2138
rect 1219 2086 1271 2138
rect 1477 2086 1529 2138
rect 1735 2086 1787 2138
rect 1993 2086 2045 2138
rect 2251 2086 2303 2138
rect 2509 2086 2561 2138
rect 2767 2086 2819 2138
rect 3025 2086 3077 2138
rect -4256 244 -3656 544
rect 6056 244 6656 544
rect 8369 85 9186 634
<< metal2 >>
rect -11156 8756 -10556 8766
rect -11156 8446 -10556 8456
rect -5444 8756 -4844 8766
rect -5444 8446 -4844 8456
rect -4256 8756 -3656 8766
rect -4256 8446 -3656 8456
rect 6056 8756 6656 8766
rect 6056 8446 6656 8456
rect 9627 7848 9867 7858
rect -3661 7671 -3393 7690
rect -3661 7468 -3641 7671
rect -3417 7468 -3393 7671
rect -3661 7450 -3393 7468
rect 7144 7642 7868 7802
rect 8028 7642 8034 7802
rect -2331 6149 645 6209
rect -2331 6097 -2245 6149
rect -2193 6097 -1987 6149
rect -1935 6097 -1729 6149
rect -1677 6097 -1471 6149
rect -1419 6097 -1213 6149
rect -1161 6097 -955 6149
rect -903 6097 -697 6149
rect -645 6097 -439 6149
rect -387 6097 -181 6149
rect -129 6097 77 6149
rect 129 6097 335 6149
rect 387 6097 593 6149
rect -2331 6089 645 6097
rect -2331 6087 926 6089
rect -2331 5991 -2235 6087
rect 525 6062 926 6087
rect 7144 6086 7304 7642
rect 9627 7595 9867 7605
rect -900 6035 -700 6045
rect -2337 5972 -2229 5991
rect -2337 5886 -2326 5972
rect -2240 5886 -2229 5972
rect -2337 5869 -2229 5886
rect 525 5916 732 6062
rect 869 5916 926 6062
rect 3600 6036 7304 6086
rect 3652 5984 5148 6036
rect 5200 5984 7304 6036
rect 3600 5926 7304 5984
rect 525 5887 926 5916
rect -900 5305 -700 5835
rect 4320 5813 4480 5823
rect 4300 5653 4320 5686
rect 4480 5653 4500 5686
rect -900 5105 700 5305
rect 500 4625 700 5105
rect 4300 4653 4500 5653
rect 500 4415 700 4425
rect 3070 4453 4500 4653
rect 3070 4376 3270 4453
rect -1232 4366 3270 4376
rect -1180 4314 -200 4366
rect -148 4314 1348 4366
rect 1400 4314 2380 4366
rect 2432 4314 3270 4366
rect -1232 4176 3270 4314
rect -1748 3048 -1696 3058
rect -1748 2148 -1696 2996
rect -716 3048 -664 3058
rect -716 2148 -664 2996
rect 316 3048 368 3058
rect 316 2148 368 2996
rect 832 3048 884 3058
rect 832 2148 884 2996
rect 1864 3048 1916 3058
rect 1864 2148 1916 2996
rect 2896 3048 2948 3058
rect 2896 2148 2948 2996
rect 3148 2450 6015 2460
rect 3388 2210 6015 2450
rect 3148 2200 6015 2210
rect -1877 2138 3077 2148
rect -1825 2086 -1619 2138
rect -1567 2086 -1361 2138
rect -1309 2086 -1103 2138
rect -1051 2086 -845 2138
rect -793 2086 -587 2138
rect -535 2086 -329 2138
rect -277 2086 -71 2138
rect -19 2086 187 2138
rect 239 2086 445 2138
rect 497 2086 703 2138
rect 755 2086 961 2138
rect 1013 2086 1219 2138
rect 1271 2086 1477 2138
rect 1529 2086 1735 2138
rect 1787 2086 1993 2138
rect 2045 2086 2251 2138
rect 2303 2086 2509 2138
rect 2561 2086 2767 2138
rect 2819 2086 3025 2138
rect -1877 2076 3077 2086
rect 5755 1536 6015 2200
rect 5755 1276 10524 1536
rect 10784 1276 10793 1536
rect 8369 634 9186 644
rect -4256 544 -3656 554
rect -4256 234 -3656 244
rect 6056 544 6656 554
rect 6056 234 6656 244
rect 8369 75 9186 85
rect -11463 -1341 -11363 -1332
rect -11728 -1363 -11628 -1354
rect -11728 -2063 -11628 -1463
rect -11732 -2153 -11723 -2063
rect -11633 -2153 -11624 -2063
rect -11463 -2085 -11363 -1441
rect -11728 -2158 -11628 -2153
rect -11467 -2175 -11458 -2085
rect -11368 -2175 -11359 -2085
rect -11463 -2180 -11363 -2175
rect -11463 -4015 -11363 -3995
rect -11463 -4095 -11453 -4015
rect -11373 -4095 -11363 -4015
rect -11713 -4826 -11633 -4816
rect -11463 -4826 -11363 -4095
rect -11633 -4906 -11363 -4826
rect -11713 -4916 -11363 -4906
<< via2 >>
rect -11156 8456 -10556 8756
rect -5444 8456 -4844 8756
rect -4256 8456 -3656 8756
rect 6056 8456 6656 8756
rect -3641 7468 -3417 7671
rect 9627 7605 9867 7848
rect -2326 5886 -2240 5972
rect 732 5916 869 6062
rect 10524 1276 10784 1536
rect -4256 244 -3656 544
rect 6056 244 6656 544
rect 8369 85 9186 634
rect -11728 -1463 -11628 -1363
rect -11463 -1441 -11363 -1341
rect -11723 -2153 -11633 -2063
rect -11458 -2175 -11368 -2085
rect -11453 -4095 -11373 -4015
rect -11713 -4906 -11633 -4826
<< metal3 >>
rect -11166 8756 -10546 8761
rect -11166 8456 -11156 8756
rect -10556 8456 -10546 8756
rect -11166 8451 -10546 8456
rect -5454 8756 -4834 8761
rect -5454 8456 -5444 8756
rect -4844 8456 -4834 8756
rect -5454 8451 -4834 8456
rect -4266 8756 -3646 8761
rect -4266 8456 -4256 8756
rect -3656 8456 -3646 8756
rect -4266 8451 -3646 8456
rect 6046 8756 6666 8761
rect 6046 8456 6056 8756
rect 6656 8456 6666 8756
rect 6046 8451 6666 8456
rect -11526 7768 -4304 8008
rect -4544 7690 -4304 7768
rect 9617 7848 9877 7853
rect -4544 7671 -3393 7690
rect -11519 7460 -11133 7560
rect -11531 7136 -11378 7236
rect -11478 1033 -11378 7136
rect -11233 1257 -11133 7460
rect -4544 7468 -3641 7671
rect -3417 7468 -3393 7671
rect 9617 7605 9627 7848
rect 9867 7840 9877 7848
rect 9867 7605 11822 7840
rect 9617 7600 11822 7605
rect -4544 7450 -3393 7468
rect 722 6062 1257 6067
rect -2337 5976 -2229 5991
rect -2337 5882 -2330 5976
rect -2236 5882 -2229 5976
rect 722 5916 732 6062
rect 869 5916 1257 6062
rect 722 5899 1257 5916
rect -2337 5869 -2229 5882
rect 1057 5312 1257 5899
rect 1057 5112 7453 5312
rect -11233 1157 -10784 1257
rect -11478 933 -10976 1033
rect -11076 -659 -10976 933
rect -11728 -759 -10976 -659
rect -11728 -1358 -11628 -759
rect -10884 -900 -10784 1157
rect -4266 544 -3646 549
rect -4266 244 -4256 544
rect -3656 244 -3646 544
rect -4266 239 -3646 244
rect 6046 544 6666 549
rect 6046 244 6056 544
rect 6656 244 6666 544
rect 6046 239 6666 244
rect 7253 -273 7453 5112
rect 10519 1536 10789 1541
rect 10519 1276 10524 1536
rect 10784 1276 11806 1536
rect 10519 1271 10789 1276
rect 8359 634 9196 639
rect 8359 85 8369 634
rect 9186 85 9196 634
rect 8359 80 9196 85
rect 7253 -473 10944 -273
rect -11463 -1000 -10784 -900
rect 10744 -714 10944 -473
rect 10744 -914 11691 -714
rect -11463 -1336 -11363 -1000
rect -11468 -1341 -11358 -1336
rect -11733 -1363 -11623 -1358
rect -11733 -1463 -11728 -1363
rect -11628 -1463 -11623 -1363
rect -11468 -1441 -11463 -1341
rect -11363 -1441 -11358 -1341
rect -11468 -1446 -11358 -1441
rect -11733 -1468 -11623 -1463
rect -11826 -1851 -11667 -1651
rect -11728 -2063 -11628 -2058
rect -11728 -2153 -11723 -2063
rect -11633 -2153 -11628 -2063
rect -11728 -4359 -11628 -2153
rect -11463 -2085 -11363 -2080
rect -11463 -2175 -11458 -2085
rect -11368 -2175 -11363 -2085
rect -11463 -4015 -11363 -2175
rect -11463 -4095 -11453 -4015
rect -11373 -4095 -11363 -4015
rect -11463 -4100 -11363 -4095
rect 11491 -4411 11691 -914
rect 11651 -4611 11691 -4411
rect -11723 -4722 -11685 -4632
rect -11723 -4826 -11623 -4722
rect -11723 -4906 -11713 -4826
rect -11633 -4906 -11623 -4826
rect -11723 -4916 -11623 -4906
<< via3 >>
rect -11156 8456 -10556 8756
rect -5444 8456 -4844 8756
rect -4256 8456 -3656 8756
rect 6056 8456 6656 8756
rect -3572 7521 -3477 7616
rect -2330 5972 -2236 5976
rect -2330 5886 -2326 5972
rect -2326 5886 -2240 5972
rect -2240 5886 -2236 5972
rect -2330 5882 -2236 5886
rect -4256 244 -3656 544
rect 6056 244 6656 544
rect 8369 85 9186 634
<< metal4 >>
rect -12000 8770 12000 9000
rect -12000 8470 -11787 8770
rect -11459 8756 12000 8770
rect -11459 8470 -11156 8756
rect -12000 8456 -11156 8470
rect -10556 8456 -5444 8756
rect -4844 8456 -4256 8756
rect -3656 8456 6056 8756
rect 6656 8456 12000 8756
rect -12000 8200 12000 8456
rect -3918 7616 -3476 7617
rect -3918 7521 -3572 7616
rect -3477 7521 -3476 7616
rect -3918 7520 -3476 7521
rect -3918 6191 -3821 7520
rect -5033 6094 -3821 6191
rect -5033 2238 -4936 6094
rect -4850 5976 -2235 5977
rect -4850 5882 -2330 5976
rect -2236 5882 -2235 5976
rect -4850 5881 -2235 5882
rect -5033 1785 -4937 2238
rect -5239 1689 -4937 1785
rect -4850 1551 -4754 5881
rect -5114 1455 -4754 1551
rect -12000 634 12000 800
rect -12000 544 8369 634
rect -12000 244 -4256 544
rect -3656 244 6056 544
rect 6656 244 8369 544
rect -12000 85 8369 244
rect 9186 85 12000 634
rect -12000 0 12000 85
<< via4 >>
rect -11787 8470 -11459 8770
rect -11756 -8756 -11428 -8456
<< metal5 >>
rect -12000 8770 -11200 9000
rect -12000 8470 -11787 8770
rect -11459 8470 -11200 8770
rect -12000 -8456 -11200 8470
rect -12000 -8756 -11756 -8456
rect -11428 -8756 -11200 -8456
rect -12000 -9000 -11200 -8756
<< comment >>
rect -850 7477 -791 7741
rect 4398 7407 4457 7671
rect 582 4226 641 4490
rect 584 2140 643 2404
use folded_cascode_n_in  folded_cascode_n_in_0 ../folded_cascode_n_in
timestamp 1622253817
transform 1 0 -3000 0 -1 -4500
box -9000 -4500 15000 4500
use sky130_fd_pr__pfet_g5v0d10v5_QFGZLW  xm4
timestamp 1621753798
transform 1 0 4400 0 1 6750
box -1901 -600 1901 600
use sky130_fd_pr__pfet_g5v0d10v5_QWKX2D  xm3
timestamp 1621753798
transform 1 0 -800 0 1 6750
box -2933 -600 2933 600
use sky130_fd_pr__nfet_g5v0d10v5_L2Y3MP  xm2
timestamp 1621753798
transform 1 0 600 0 1 1500
box -2867 -588 2867 588
use sky130_fd_pr__nfet_g5v0d10v5_DQEKTK  xm1
timestamp 1621753798
transform 1 0 600 0 1 3600
box -3899 -588 3899 588
use sky130_fd_pr__res_high_po_1p41_30um  sky130_fd_pr__res_high_po_1p41_30um_2
timestamp 1621758535
transform 1 0 9400 0 1 4500
box -143 -3432 143 3432
use sky130_fd_pr__res_high_po_1p41_30um  sky130_fd_pr__res_high_po_1p41_30um_1
timestamp 1621758535
transform 1 0 8800 0 1 4500
box -143 -3432 143 3432
use sky130_fd_pr__res_high_po_1p41_30um  sky130_fd_pr__res_high_po_1p41_30um_0
timestamp 1621758535
transform 1 0 8200 0 1 4500
box -143 -3432 143 3432
use sky130_fd_pr__cap_mim_m3_1_28umx28um  sky130_fd_pr__cap_mim_m3_1_28umx28um_0
timestamp 1621745012
transform 0 1 -8050 -1 0 4450
box -3000 -2950 2999 2950
<< labels >>
flabel metal4 -12000 8200 -12000 9000 3 FreeSans 480 0 0 0 vdd
port 7 e
flabel metal4 -12000 0 -12000 800 3 FreeSans 480 0 0 0 vss
port 8 e
flabel metal3 11806 1276 11806 1536 1 FreeSans 240 0 0 0 imon
port 2 n
flabel metal3 11822 7600 11822 7840 1 FreeSans 240 0 0 0 isense
port 3 n
flabel metal3 -11826 -1851 -11826 -1651 0 FreeSans 240 0 0 0 ibias
port 1 nsew
flabel metal3 s -11526 7768 -11523 8008 0 FreeSans 240 0 0 0 sense_fet
port 4 nsew
flabel metal3 s -11519 7460 -11517 7560 0 FreeSans 240 0 0 0 sense_fet_kelvin
port 5 nsew
flabel metal3 s -11531 7136 -11526 7236 0 FreeSans 240 0 0 0 sw_node
port 6 nsew
<< properties >>
string FIXED_BBOX -11242 1158 -4758 8842
<< end >>
