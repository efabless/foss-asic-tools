magic
tech sky130A
magscale 1 2
timestamp 1621739502
<< nwell >>
rect -3000 40 3000 4500
<< pwell >>
rect -3000 -4500 3000 -40
<< mvpsubdiff >>
rect -2934 -118 2934 -106
rect -2934 -278 -2700 -118
rect 2700 -278 2934 -118
rect -2934 -290 2934 -278
rect -2934 -340 -2750 -290
rect -2934 -4200 -2922 -340
rect -2762 -4200 -2750 -340
rect -2934 -4250 -2750 -4200
rect 2750 -340 2934 -290
rect 2750 -4200 2762 -340
rect 2922 -4200 2934 -340
rect 2750 -4250 2934 -4200
rect -2934 -4262 2934 -4250
rect -2934 -4422 -2700 -4262
rect 2700 -4422 2934 -4262
rect -2934 -4434 2934 -4422
<< mvnsubdiff >>
rect -2934 4422 2934 4434
rect -2934 4262 -2700 4422
rect 2700 4262 2934 4422
rect -2934 4250 2934 4262
rect -2934 4200 -2750 4250
rect -2934 340 -2922 4200
rect -2762 340 -2750 4200
rect -2934 290 -2750 340
rect 2750 4200 2934 4250
rect 2750 340 2762 4200
rect 2922 340 2934 4200
rect 2750 290 2934 340
rect -2934 278 2934 290
rect -2934 118 -2700 278
rect 2700 118 2934 278
rect -2934 106 2934 118
<< mvpsubdiffcont >>
rect -2700 -278 2700 -118
rect -2922 -4200 -2762 -340
rect 2762 -4200 2922 -340
rect -2700 -4422 2700 -4262
<< mvnsubdiffcont >>
rect -2700 4262 2700 4422
rect -2922 340 -2762 4200
rect 2762 340 2922 4200
rect -2700 118 2700 278
<< locali >>
rect -2922 4200 -2762 4422
rect 2762 4200 2922 4422
rect -1227 1259 1227 1453
rect -2922 118 -2762 340
rect 2762 118 2922 340
rect -2922 -340 -2762 -118
rect 2762 -340 2922 -118
rect -2259 -1462 2259 -1107
rect -2922 -4422 -2762 -4200
rect 2762 -4422 2922 -4200
<< viali >>
rect -2762 4262 -2700 4422
rect -2700 4262 2700 4422
rect 2700 4262 2762 4422
rect -2922 477 -2762 4063
rect 2762 477 2922 4063
rect -2762 118 -2700 278
rect -2700 118 2700 278
rect 2700 118 2762 278
rect -2762 -278 -2700 -118
rect -2700 -278 2700 -118
rect 2700 -278 2762 -118
rect -2922 -4063 -2762 -477
rect 2762 -4063 2922 -477
rect -2762 -4422 -2700 -4262
rect -2700 -4422 2700 -4262
rect 2700 -4422 2762 -4262
<< metal1 >>
rect -2928 4422 2928 4428
rect -2928 4262 -2762 4422
rect 2762 4262 2928 4422
rect -2928 4256 2928 4262
rect -2928 4063 -2756 4256
rect -2928 477 -2922 4063
rect -2762 3956 -2756 4063
rect -2156 3956 2156 4256
rect 2756 4063 2928 4256
rect 2756 3956 2762 4063
rect -2762 2866 2762 3956
rect -2762 477 -2756 2866
rect -1571 2587 -1525 2866
rect -1313 2587 -1267 2866
rect -1571 2541 -1267 2587
rect -1571 2500 -1525 2541
rect -1313 2500 -1267 2541
rect -797 2500 -751 2866
rect -281 2500 -235 2866
rect 235 2500 281 2866
rect 751 2500 797 2866
rect 1267 2587 1313 2866
rect 1525 2587 1571 2866
rect 1267 2541 1571 2587
rect 1267 2500 1313 2541
rect 1525 2500 1571 2541
rect -1055 1130 -1009 1500
rect -539 1330 -493 1500
rect -23 1459 23 1500
rect -175 1413 175 1459
rect -556 1270 -546 1330
rect -486 1270 -476 1330
rect -1072 1070 -1062 1130
rect -1002 1070 -992 1130
rect -23 930 23 1413
rect 493 1130 539 1500
rect 1009 1330 1055 1500
rect 992 1270 1002 1330
rect 1062 1270 1072 1330
rect 476 1070 486 1130
rect 546 1070 556 1130
rect -60 830 -50 930
rect 50 830 60 930
rect -2928 284 -2756 477
rect 2756 477 2762 2866
rect 2922 477 2928 4063
rect 2756 284 2928 477
rect -2928 278 2928 284
rect -2928 118 -2762 278
rect 2762 118 2928 278
rect -2928 112 2928 118
rect -2928 -118 2928 -112
rect -2928 -278 -2762 -118
rect 2762 -278 2928 -118
rect -2928 -284 2928 -278
rect -2928 -477 -2756 -284
rect -2928 -4063 -2922 -477
rect -2762 -2822 -2756 -477
rect 2756 -477 2928 -284
rect -60 -860 -50 -760
rect 50 -860 60 -760
rect -576 -1010 -566 -910
rect -466 -1010 -456 -910
rect -539 -1500 -493 -1010
rect -23 -1500 23 -860
rect 972 -1180 982 -1080
rect 1082 -1180 1092 -1080
rect 456 -1350 466 -1250
rect 566 -1350 576 -1250
rect 493 -1500 539 -1350
rect 1009 -1500 1055 -1180
rect -2603 -2532 -2557 -2500
rect -2345 -2532 -2299 -2500
rect -2087 -2532 -2041 -2500
rect -2603 -2634 -2299 -2532
rect -2239 -2578 -1889 -2532
rect -2603 -2822 -2557 -2634
rect -2345 -2822 -2299 -2634
rect -2087 -2670 -2041 -2578
rect -2104 -2730 -2094 -2670
rect -2034 -2730 -2024 -2670
rect -1829 -2822 -1783 -2500
rect -1571 -2532 -1525 -2500
rect -1723 -2578 -1373 -2532
rect -1571 -2670 -1525 -2578
rect -1588 -2730 -1578 -2670
rect -1518 -2730 -1508 -2670
rect -1313 -2822 -1267 -2500
rect -1055 -2532 -1009 -2500
rect -1207 -2578 -857 -2532
rect -1055 -2670 -1009 -2578
rect -1072 -2730 -1062 -2670
rect -1002 -2730 -992 -2670
rect -797 -2822 -751 -2500
rect -281 -2822 -235 -2500
rect 235 -2822 281 -2500
rect 751 -2822 797 -2500
rect 1267 -2822 1313 -2500
rect 1525 -2532 1571 -2500
rect 1373 -2578 1723 -2532
rect 1525 -2670 1571 -2578
rect 1508 -2730 1518 -2670
rect 1578 -2730 1588 -2670
rect 1783 -2822 1829 -2500
rect 2041 -2532 2087 -2500
rect 2299 -2532 2345 -2500
rect 2557 -2532 2603 -2500
rect 1889 -2578 2239 -2532
rect 2041 -2670 2087 -2578
rect 2299 -2637 2603 -2532
rect 2024 -2730 2034 -2670
rect 2094 -2730 2104 -2670
rect 2299 -2822 2345 -2637
rect 2557 -2822 2603 -2637
rect 2756 -2822 2762 -477
rect -2762 -3956 2762 -2822
rect -2762 -4063 -2756 -3956
rect -2928 -4256 -2756 -4063
rect -2156 -4256 2156 -3956
rect 2756 -4063 2762 -3956
rect 2922 -4063 2928 -477
rect 2756 -4256 2928 -4063
rect -2928 -4262 2928 -4256
rect -2928 -4422 -2762 -4262
rect 2762 -4422 2928 -4262
rect -2928 -4428 2928 -4422
<< via1 >>
rect -2756 3956 -2156 4256
rect 2156 3956 2756 4256
rect -546 1270 -486 1330
rect -1062 1070 -1002 1130
rect 1002 1270 1062 1330
rect 486 1070 546 1130
rect -50 830 50 930
rect -50 -860 50 -760
rect -566 -1010 -466 -910
rect 982 -1180 1082 -1080
rect 466 -1350 566 -1250
rect -2094 -2730 -2034 -2670
rect -1578 -2730 -1518 -2670
rect -1062 -2730 -1002 -2670
rect 1518 -2730 1578 -2670
rect 2034 -2730 2094 -2670
rect -2756 -4256 -2156 -3956
rect 2156 -4256 2756 -3956
<< metal2 >>
rect -2756 4256 -2156 4266
rect -2756 3946 -2156 3956
rect 2156 4256 2756 4266
rect 2156 3946 2756 3956
rect 962 1340 1062 1350
rect -546 1330 962 1340
rect -486 1270 962 1330
rect -546 1260 962 1270
rect 962 1230 1062 1240
rect 446 1140 546 1150
rect -1062 1130 446 1140
rect -1002 1070 446 1130
rect -1062 1060 446 1070
rect 446 1030 546 1040
rect -50 930 50 940
rect -50 -760 50 830
rect -50 -870 50 -860
rect -566 -910 -466 -900
rect -566 -1020 -466 -1010
rect 982 -1080 1082 -1070
rect 982 -1190 1082 -1180
rect 466 -1250 566 -1240
rect 466 -1360 566 -1350
rect -2094 -2670 2094 -2660
rect -2034 -2730 -1578 -2670
rect -1518 -2730 -1062 -2670
rect -1002 -2730 1518 -2670
rect 1578 -2730 2034 -2670
rect -2094 -2780 2094 -2730
rect -2094 -2960 -100 -2780
rect 100 -2960 2094 -2780
rect -100 -2990 100 -2980
rect -2756 -3956 -2156 -3946
rect -2756 -4266 -2156 -4256
rect 2156 -3956 2756 -3946
rect 2156 -4266 2756 -4256
<< via2 >>
rect -2756 3956 -2156 4256
rect 2156 3956 2756 4256
rect 962 1330 1062 1340
rect 962 1270 1002 1330
rect 1002 1270 1062 1330
rect 962 1240 1062 1270
rect 446 1130 546 1140
rect 446 1070 486 1130
rect 486 1070 546 1130
rect 446 1040 546 1070
rect -566 -1010 -466 -910
rect 982 -1180 1082 -1080
rect 466 -1350 566 -1250
rect -100 -2980 100 -2780
rect -2756 -4256 -2156 -3956
rect 2156 -4256 2756 -3956
<< metal3 >>
rect -2766 4256 -2146 4261
rect -2766 3956 -2756 4256
rect -2156 3956 -2146 4256
rect -2766 3951 -2146 3956
rect 2146 4256 2766 4261
rect 2146 3956 2156 4256
rect 2756 3956 2766 4256
rect 2146 3951 2766 3956
rect 952 1340 1908 1345
rect 952 1240 962 1340
rect 1062 1240 1908 1340
rect 952 1235 1908 1240
rect 436 1140 1911 1145
rect 436 1040 446 1140
rect 546 1040 1911 1140
rect 436 1035 1911 1040
rect -576 -910 -456 -905
rect -576 -1010 -566 -910
rect -466 -1010 2446 -910
rect -576 -1015 -456 -1010
rect 972 -1080 1092 -1075
rect 972 -1180 982 -1080
rect 1082 -1180 2449 -1080
rect 972 -1185 1092 -1180
rect 456 -1250 576 -1245
rect 456 -1350 466 -1250
rect 566 -1350 2449 -1250
rect 456 -1355 576 -1350
rect -110 -2780 110 -2775
rect -2528 -2980 -100 -2780
rect 100 -2980 110 -2780
rect -110 -2985 110 -2980
rect -2766 -3956 -2146 -3951
rect -2766 -4256 -2756 -3956
rect -2156 -4256 -2146 -3956
rect -2766 -4261 -2146 -4256
rect 2146 -3956 2766 -3951
rect 2146 -4256 2156 -3956
rect 2756 -4256 2766 -3956
rect 2146 -4261 2766 -4256
<< via3 >>
rect -2756 3956 -2156 4256
rect 2156 3956 2756 4256
rect -2756 -4256 -2156 -3956
rect 2156 -4256 2756 -3956
<< metal4 >>
rect -3000 4256 3000 4500
rect -3000 3956 -2756 4256
rect -2156 3956 2156 4256
rect 2756 3956 3000 4256
rect -3000 3700 3000 3956
rect -3000 -3956 3000 -3700
rect -3000 -4256 -2756 -3956
rect -2156 -4256 2156 -3956
rect 2756 -4256 3000 -3956
rect -3000 -4500 3000 -4256
use sky130_fd_pr__pfet_g5v0d10v5_QNH2MW  xm2
timestamp 1621737489
transform 1 0 0 0 1 2000
box -1643 -600 1643 600
use sky130_fd_pr__nfet_g5v0d10v5_DQEKPQ  xm1
timestamp 1621737489
transform 1 0 0 0 1 -2000
box -2609 -588 2609 588
<< labels >>
flabel metal4 -3000 3700 -3000 4500 3 FreeSans 480 0 0 0 vdd
port 7 e
flabel metal4 -3000 -4500 -3000 -3700 3 FreeSans 480 0 0 0 vss
port 8 e
flabel metal3 1908 1235 1908 1345 1 FreeSans 240 0 0 0 bias_opa_n
port 5 n
flabel metal3 1911 1035 1911 1145 1 FreeSans 240 0 0 0 bias_opa_p
port 6 n
flabel metal3 2446 -1010 2446 -910 1 FreeSans 240 0 0 0 bias_current_shift
port 3 n
flabel metal3 2449 -1180 2449 -1080 1 FreeSans 240 0 0 0 bias_cmp_2
port 2 n
flabel metal3 2449 -1350 2449 -1250 1 FreeSans 240 0 0 0 bias_cmp
port 1 n
flabel metal3 -2528 -2980 -2528 -2780 1 FreeSans 240 0 0 0 bias_in
port 4 n
<< properties >>
string FIXED_BBOX -2842 -4342 2842 -198
<< end >>
