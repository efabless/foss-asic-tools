MACRO INVERTER
  ORIGIN 0 0 ;
  FOREIGN INVERTER 0 0 ;
  SIZE 13.02 BY 14.03 ;
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 0.26 3.58 6.46 ;
      LAYER M3 ;
        RECT 8.46 0.26 8.74 6.46 ;
      LAYER M3 ;
        RECT 3.3 1.075 3.58 1.445 ;
      LAYER M2 ;
        RECT 3.44 1.12 8.6 1.4 ;
      LAYER M3 ;
        RECT 8.46 1.075 8.74 1.445 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 2.87 4.46 3.15 10.66 ;
      LAYER M3 ;
        RECT 8.89 4.46 9.17 10.66 ;
      LAYER M3 ;
        RECT 2.87 4.855 3.15 5.225 ;
      LAYER M2 ;
        RECT 3.01 4.9 9.03 5.18 ;
      LAYER M3 ;
        RECT 8.89 4.855 9.17 5.225 ;
    END
  END A
  OBS 
  LAYER M1 ;
        RECT 7.185 0.335 7.435 3.865 ;
  LAYER M1 ;
        RECT 7.185 4.115 7.435 5.125 ;
  LAYER M1 ;
        RECT 7.185 6.215 7.435 9.745 ;
  LAYER M1 ;
        RECT 7.185 9.995 7.435 11.005 ;
  LAYER M1 ;
        RECT 7.185 12.095 7.435 13.105 ;
  LAYER M1 ;
        RECT 6.755 0.335 7.005 3.865 ;
  LAYER M1 ;
        RECT 6.755 6.215 7.005 9.745 ;
  LAYER M1 ;
        RECT 7.615 0.335 7.865 3.865 ;
  LAYER M1 ;
        RECT 7.615 6.215 7.865 9.745 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 3.865 ;
  LAYER M1 ;
        RECT 8.045 4.115 8.295 5.125 ;
  LAYER M1 ;
        RECT 8.045 6.215 8.295 9.745 ;
  LAYER M1 ;
        RECT 8.045 9.995 8.295 11.005 ;
  LAYER M1 ;
        RECT 8.045 12.095 8.295 13.105 ;
  LAYER M1 ;
        RECT 8.475 0.335 8.725 3.865 ;
  LAYER M1 ;
        RECT 8.475 6.215 8.725 9.745 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 3.865 ;
  LAYER M1 ;
        RECT 8.905 4.115 9.155 5.125 ;
  LAYER M1 ;
        RECT 8.905 6.215 9.155 9.745 ;
  LAYER M1 ;
        RECT 8.905 9.995 9.155 11.005 ;
  LAYER M1 ;
        RECT 8.905 12.095 9.155 13.105 ;
  LAYER M1 ;
        RECT 9.335 0.335 9.585 3.865 ;
  LAYER M1 ;
        RECT 9.335 6.215 9.585 9.745 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 3.865 ;
  LAYER M1 ;
        RECT 9.765 4.115 10.015 5.125 ;
  LAYER M1 ;
        RECT 9.765 6.215 10.015 9.745 ;
  LAYER M1 ;
        RECT 9.765 9.995 10.015 11.005 ;
  LAYER M1 ;
        RECT 9.765 12.095 10.015 13.105 ;
  LAYER M1 ;
        RECT 10.195 0.335 10.445 3.865 ;
  LAYER M1 ;
        RECT 10.195 6.215 10.445 9.745 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 3.865 ;
  LAYER M1 ;
        RECT 10.625 4.115 10.875 5.125 ;
  LAYER M1 ;
        RECT 10.625 6.215 10.875 9.745 ;
  LAYER M1 ;
        RECT 10.625 9.995 10.875 11.005 ;
  LAYER M1 ;
        RECT 10.625 12.095 10.875 13.105 ;
  LAYER M1 ;
        RECT 11.055 0.335 11.305 3.865 ;
  LAYER M1 ;
        RECT 11.055 6.215 11.305 9.745 ;
  LAYER M2 ;
        RECT 7.14 0.28 10.92 0.56 ;
  LAYER M2 ;
        RECT 7.14 4.48 10.92 4.76 ;
  LAYER M2 ;
        RECT 6.71 0.7 11.35 0.98 ;
  LAYER M2 ;
        RECT 7.14 6.16 10.92 6.44 ;
  LAYER M2 ;
        RECT 7.14 10.36 10.92 10.64 ;
  LAYER M2 ;
        RECT 7.14 12.46 10.92 12.74 ;
  LAYER M2 ;
        RECT 6.71 6.58 11.35 6.86 ;
  LAYER M3 ;
        RECT 8.46 0.26 8.74 6.46 ;
  LAYER M3 ;
        RECT 8.89 4.46 9.17 10.66 ;
  LAYER M3 ;
        RECT 9.32 0.68 9.6 12.76 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 3.865 ;
  LAYER M1 ;
        RECT 4.605 4.115 4.855 5.125 ;
  LAYER M1 ;
        RECT 4.605 6.215 4.855 9.745 ;
  LAYER M1 ;
        RECT 4.605 9.995 4.855 11.005 ;
  LAYER M1 ;
        RECT 4.605 12.095 4.855 13.105 ;
  LAYER M1 ;
        RECT 5.035 0.335 5.285 3.865 ;
  LAYER M1 ;
        RECT 5.035 6.215 5.285 9.745 ;
  LAYER M1 ;
        RECT 4.175 0.335 4.425 3.865 ;
  LAYER M1 ;
        RECT 4.175 6.215 4.425 9.745 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 3.865 ;
  LAYER M1 ;
        RECT 3.745 4.115 3.995 5.125 ;
  LAYER M1 ;
        RECT 3.745 6.215 3.995 9.745 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 12.095 3.995 13.105 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 3.865 ;
  LAYER M1 ;
        RECT 3.315 6.215 3.565 9.745 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 3.865 ;
  LAYER M1 ;
        RECT 2.885 4.115 3.135 5.125 ;
  LAYER M1 ;
        RECT 2.885 6.215 3.135 9.745 ;
  LAYER M1 ;
        RECT 2.885 9.995 3.135 11.005 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 13.105 ;
  LAYER M1 ;
        RECT 2.455 0.335 2.705 3.865 ;
  LAYER M1 ;
        RECT 2.455 6.215 2.705 9.745 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 3.865 ;
  LAYER M1 ;
        RECT 2.025 4.115 2.275 5.125 ;
  LAYER M1 ;
        RECT 2.025 6.215 2.275 9.745 ;
  LAYER M1 ;
        RECT 2.025 9.995 2.275 11.005 ;
  LAYER M1 ;
        RECT 2.025 12.095 2.275 13.105 ;
  LAYER M1 ;
        RECT 1.595 0.335 1.845 3.865 ;
  LAYER M1 ;
        RECT 1.595 6.215 1.845 9.745 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 3.865 ;
  LAYER M1 ;
        RECT 1.165 4.115 1.415 5.125 ;
  LAYER M1 ;
        RECT 1.165 6.215 1.415 9.745 ;
  LAYER M1 ;
        RECT 1.165 9.995 1.415 11.005 ;
  LAYER M1 ;
        RECT 1.165 12.095 1.415 13.105 ;
  LAYER M1 ;
        RECT 0.735 0.335 0.985 3.865 ;
  LAYER M1 ;
        RECT 0.735 6.215 0.985 9.745 ;
  LAYER M2 ;
        RECT 1.12 0.28 4.9 0.56 ;
  LAYER M2 ;
        RECT 1.12 4.48 4.9 4.76 ;
  LAYER M2 ;
        RECT 0.69 0.7 5.33 0.98 ;
  LAYER M2 ;
        RECT 1.12 6.16 4.9 6.44 ;
  LAYER M2 ;
        RECT 1.12 10.36 4.9 10.64 ;
  LAYER M2 ;
        RECT 1.12 12.46 4.9 12.74 ;
  LAYER M2 ;
        RECT 0.69 6.58 5.33 6.86 ;
  LAYER M3 ;
        RECT 3.3 0.26 3.58 6.46 ;
  LAYER M3 ;
        RECT 2.87 4.46 3.15 10.66 ;
  LAYER M3 ;
        RECT 2.44 0.68 2.72 12.76 ;
  END 
END INVERTER
