** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom8k.sch
**.subckt rom8k
*+ LDQ[15],LDQ[14],LDQ[13],LDQ[12],LDQ[11],LDQ[10],LDQ[9],LDQ[8],LDQ[7],LDQ[6],LDQ[5],LDQ[4],LDQ[3],LDQ[2],LDQ[1],LDQ[0] LDA[12],LDA[11],LDA[10],LDA[9],LDA[8],LDA[7],LDA[6],LDA[5],LDA[4],LDA[3],LDA[2],LDA[1],LDA[0] LDCP
*+ LDEN LDOE vss vcc
*.opin
*+ LDQ[15],LDQ[14],LDQ[13],LDQ[12],LDQ[11],LDQ[10],LDQ[9],LDQ[8],LDQ[7],LDQ[6],LDQ[5],LDQ[4],LDQ[3],LDQ[2],LDQ[1],LDQ[0]
*.ipin LDA[12],LDA[11],LDA[10],LDA[9],LDA[8],LDA[7],LDA[6],LDA[5],LDA[4],LDA[3],LDA[2],LDA[1],LDA[0]
*.ipin LDCP
*.ipin LDEN
*.ipin LDOE
*.ipin vss
*.ipin vcc
xcdec[15] LDYMS[15] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[255] LDBL[254] LDBL[253] LDBL[252] LDBL[251]
+ LDBL[250] LDBL[249] LDBL[248] LDBL[247] LDBL[246] LDBL[245] LDBL[244] LDBL[243] LDBL[242] LDBL[241] LDBL[240]
+ vss rom2_coldec
xcdec[14] LDYMS[14] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[239] LDBL[238] LDBL[237] LDBL[236] LDBL[235]
+ LDBL[234] LDBL[233] LDBL[232] LDBL[231] LDBL[230] LDBL[229] LDBL[228] LDBL[227] LDBL[226] LDBL[225] LDBL[224]
+ vss rom2_coldec
xcdec[13] LDYMS[13] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[223] LDBL[222] LDBL[221] LDBL[220] LDBL[219]
+ LDBL[218] LDBL[217] LDBL[216] LDBL[215] LDBL[214] LDBL[213] LDBL[212] LDBL[211] LDBL[210] LDBL[209] LDBL[208]
+ vss rom2_coldec
xcdec[12] LDYMS[12] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[207] LDBL[206] LDBL[205] LDBL[204] LDBL[203]
+ LDBL[202] LDBL[201] LDBL[200] LDBL[199] LDBL[198] LDBL[197] LDBL[196] LDBL[195] LDBL[194] LDBL[193] LDBL[192]
+ vss rom2_coldec
xcdec[11] LDYMS[11] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[191] LDBL[190] LDBL[189] LDBL[188] LDBL[187]
+ LDBL[186] LDBL[185] LDBL[184] LDBL[183] LDBL[182] LDBL[181] LDBL[180] LDBL[179] LDBL[178] LDBL[177] LDBL[176]
+ vss rom2_coldec
xcdec[10] LDYMS[10] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[175] LDBL[174] LDBL[173] LDBL[172] LDBL[171]
+ LDBL[170] LDBL[169] LDBL[168] LDBL[167] LDBL[166] LDBL[165] LDBL[164] LDBL[163] LDBL[162] LDBL[161] LDBL[160]
+ vss rom2_coldec
xcdec[9] LDYMS[9] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[159] LDBL[158] LDBL[157] LDBL[156] LDBL[155]
+ LDBL[154] LDBL[153] LDBL[152] LDBL[151] LDBL[150] LDBL[149] LDBL[148] LDBL[147] LDBL[146] LDBL[145] LDBL[144]
+ vss rom2_coldec
xcdec[8] LDYMS[8] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[143] LDBL[142] LDBL[141] LDBL[140] LDBL[139]
+ LDBL[138] LDBL[137] LDBL[136] LDBL[135] LDBL[134] LDBL[133] LDBL[132] LDBL[131] LDBL[130] LDBL[129] LDBL[128]
+ vss rom2_coldec
xcdec[7] LDYMS[7] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[127] LDBL[126] LDBL[125] LDBL[124] LDBL[123]
+ LDBL[122] LDBL[121] LDBL[120] LDBL[119] LDBL[118] LDBL[117] LDBL[116] LDBL[115] LDBL[114] LDBL[113] LDBL[112]
+ vss rom2_coldec
xcdec[6] LDYMS[6] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[111] LDBL[110] LDBL[109] LDBL[108] LDBL[107]
+ LDBL[106] LDBL[105] LDBL[104] LDBL[103] LDBL[102] LDBL[101] LDBL[100] LDBL[99] LDBL[98] LDBL[97] LDBL[96] vss
+ rom2_coldec
xcdec[5] LDYMS[5] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[95] LDBL[94] LDBL[93] LDBL[92] LDBL[91]
+ LDBL[90] LDBL[89] LDBL[88] LDBL[87] LDBL[86] LDBL[85] LDBL[84] LDBL[83] LDBL[82] LDBL[81] LDBL[80] vss
+ rom2_coldec
xcdec[4] LDYMS[4] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[79] LDBL[78] LDBL[77] LDBL[76] LDBL[75]
+ LDBL[74] LDBL[73] LDBL[72] LDBL[71] LDBL[70] LDBL[69] LDBL[68] LDBL[67] LDBL[66] LDBL[65] LDBL[64] vss
+ rom2_coldec
xcdec[3] LDYMS[3] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[63] LDBL[62] LDBL[61] LDBL[60] LDBL[59]
+ LDBL[58] LDBL[57] LDBL[56] LDBL[55] LDBL[54] LDBL[53] LDBL[52] LDBL[51] LDBL[50] LDBL[49] LDBL[48] vss
+ rom2_coldec
xcdec[2] LDYMS[2] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[47] LDBL[46] LDBL[45] LDBL[44] LDBL[43]
+ LDBL[42] LDBL[41] LDBL[40] LDBL[39] LDBL[38] LDBL[37] LDBL[36] LDBL[35] LDBL[34] LDBL[33] LDBL[32] vss
+ rom2_coldec
xcdec[1] LDYMS[1] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[31] LDBL[30] LDBL[29] LDBL[28] LDBL[27]
+ LDBL[26] LDBL[25] LDBL[24] LDBL[23] LDBL[22] LDBL[21] LDBL[20] LDBL[19] LDBL[18] LDBL[17] LDBL[16] vss
+ rom2_coldec
xcdec[0] LDYMS[0] LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7]
+ LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[15] LDBL[14] LDBL[13] LDBL[12] LDBL[11]
+ LDBL[10] LDBL[9] LDBL[8] LDBL[7] LDBL[6] LDBL[5] LDBL[4] LDBL[3] LDBL[2] LDBL[1] LDBL[0] vss rom2_coldec
xsa[15] LDQ[15] LDCP_SA LDYMS[15] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[14] LDQ[14] LDCP_SA LDYMS[14] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[13] LDQ[13] LDCP_SA LDYMS[13] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[12] LDQ[12] LDCP_SA LDYMS[12] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[11] LDQ[11] LDCP_SA LDYMS[11] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[10] LDQ[10] LDCP_SA LDYMS[10] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[9] LDQ[9] LDCP_SA LDYMS[9] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[8] LDQ[8] LDCP_SA LDYMS[8] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[7] LDQ[7] LDCP_SA LDYMS[7] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[6] LDQ[6] LDCP_SA LDYMS[6] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[5] LDQ[5] LDCP_SA LDYMS[5] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[4] LDQ[4] LDCP_SA LDYMS[4] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[3] LDQ[3] LDCP_SA LDYMS[3] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[2] LDQ[2] LDCP_SA LDYMS[2] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[1] LDQ[1] LDCP_SA LDYMS[1] LDOE LDPRECH LDSAL vccsa vss rom2_sa
xsa[0] LDQ[0] LDCP_SA LDYMS[0] LDOE LDPRECH LDSAL vccsa vss rom2_sa
vsa vcc vccsa 0
vdec vcc vccdec 0
vl vcc vccl 0
xlat LDEN_LAT LDAI[12] LDAI[11] LDAI[10] LDAI[9] LDAI[8] LDAI[7] LDAI[6] LDAI[5] LDAI[4] LDAI[3]
+ LDAI[2] LDAI[1] LDAI[0] LDEN LDCP_ADDLAT_B LDA[12] LDA[11] LDA[10] LDA[9] LDA[8] LDA[7] LDA[6] LDA[5]
+ LDA[4] LDA[3] LDA[2] LDA[1] LDA[0] vccl vss rom2_addlatch
xctrl LDPRECH LDSAL LDCP_ROWDEC LDCP_SA LDCP_ADDLAT_B LDCP_COL_B LDEN_LAT LDCP vccl vss LDYMSREF
+ rom2_ctrl
xcpre LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8] LDY1[7] LDY1[6] LDY1[5]
+ LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDAI[3] LDAI[2] LDAI[1] LDAI[0] vccdec vss rom2_predec3
c1[15] LDL1X[15] vss 210f m=1
c1[14] LDL1X[14] vss 210f m=1
c1[13] LDL1X[13] vss 210f m=1
c1[12] LDL1X[12] vss 210f m=1
c1[11] LDL1X[11] vss 210f m=1
c1[10] LDL1X[10] vss 210f m=1
c1[9] LDL1X[9] vss 210f m=1
c1[8] LDL1X[8] vss 210f m=1
c1[7] LDL1X[7] vss 210f m=1
c1[6] LDL1X[6] vss 210f m=1
c1[5] LDL1X[5] vss 210f m=1
c1[4] LDL1X[4] vss 210f m=1
c1[3] LDL1X[3] vss 210f m=1
c1[2] LDL1X[2] vss 210f m=1
c1[1] LDL1X[1] vss 210f m=1
c1[0] LDL1X[0] vss 210f m=1
c2[3] LDL2X[3] vss 120f m=1
c2[2] LDL2X[2] vss 120f m=1
c2[1] LDL2X[1] vss 120f m=1
c2[0] LDL2X[0] vss 120f m=1
c4[12] LDAI[12] vss 40f m=1
c4[11] LDAI[11] vss 40f m=1
c4[10] LDAI[10] vss 40f m=1
c4[9] LDAI[9] vss 40f m=1
c4[8] LDAI[8] vss 40f m=1
c4[7] LDAI[7] vss 40f m=1
c4[6] LDAI[6] vss 40f m=1
c4[5] LDAI[5] vss 40f m=1
c4[4] LDAI[4] vss 40f m=1
c4[3] LDAI[3] vss 40f m=1
c4[2] LDAI[2] vss 40f m=1
c4[1] LDAI[1] vss 40f m=1
c4[0] LDAI[0] vss 40f m=1
c5[15] LDY1[15] vss 45f m=1
c5[14] LDY1[14] vss 45f m=1
c5[13] LDY1[13] vss 45f m=1
c5[12] LDY1[12] vss 45f m=1
c5[11] LDY1[11] vss 45f m=1
c5[10] LDY1[10] vss 45f m=1
c5[9] LDY1[9] vss 45f m=1
c5[8] LDY1[8] vss 45f m=1
c5[7] LDY1[7] vss 45f m=1
c5[6] LDY1[6] vss 45f m=1
c5[5] LDY1[5] vss 45f m=1
c5[4] LDY1[4] vss 45f m=1
c5[3] LDY1[3] vss 45f m=1
c5[2] LDY1[2] vss 45f m=1
c5[1] LDY1[1] vss 45f m=1
c5[0] LDY1[0] vss 45f m=1
xrdec[31] LDWL[511] LDWL[510] LDWL[509] LDWL[508] LDWL[507] LDWL[506] LDWL[505] LDWL[504] LDWL[503]
+ LDWL[502] LDWL[501] LDWL[500] LDWL[499] LDWL[498] LDWL[497] LDWL[496] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[3] LDL3X[7] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[30] LDWL[495] LDWL[494] LDWL[493] LDWL[492] LDWL[491] LDWL[490] LDWL[489] LDWL[488] LDWL[487]
+ LDWL[486] LDWL[485] LDWL[484] LDWL[483] LDWL[482] LDWL[481] LDWL[480] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[2] LDL3X[7] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[29] LDWL[479] LDWL[478] LDWL[477] LDWL[476] LDWL[475] LDWL[474] LDWL[473] LDWL[472] LDWL[471]
+ LDWL[470] LDWL[469] LDWL[468] LDWL[467] LDWL[466] LDWL[465] LDWL[464] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[1] LDL3X[7] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[28] LDWL[463] LDWL[462] LDWL[461] LDWL[460] LDWL[459] LDWL[458] LDWL[457] LDWL[456] LDWL[455]
+ LDWL[454] LDWL[453] LDWL[452] LDWL[451] LDWL[450] LDWL[449] LDWL[448] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[0] LDL3X[7] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[27] LDWL[447] LDWL[446] LDWL[445] LDWL[444] LDWL[443] LDWL[442] LDWL[441] LDWL[440] LDWL[439]
+ LDWL[438] LDWL[437] LDWL[436] LDWL[435] LDWL[434] LDWL[433] LDWL[432] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[3] LDL3X[6] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[26] LDWL[431] LDWL[430] LDWL[429] LDWL[428] LDWL[427] LDWL[426] LDWL[425] LDWL[424] LDWL[423]
+ LDWL[422] LDWL[421] LDWL[420] LDWL[419] LDWL[418] LDWL[417] LDWL[416] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[2] LDL3X[6] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[25] LDWL[415] LDWL[414] LDWL[413] LDWL[412] LDWL[411] LDWL[410] LDWL[409] LDWL[408] LDWL[407]
+ LDWL[406] LDWL[405] LDWL[404] LDWL[403] LDWL[402] LDWL[401] LDWL[400] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[1] LDL3X[6] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[24] LDWL[399] LDWL[398] LDWL[397] LDWL[396] LDWL[395] LDWL[394] LDWL[393] LDWL[392] LDWL[391]
+ LDWL[390] LDWL[389] LDWL[388] LDWL[387] LDWL[386] LDWL[385] LDWL[384] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[0] LDL3X[6] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[23] LDWL[383] LDWL[382] LDWL[381] LDWL[380] LDWL[379] LDWL[378] LDWL[377] LDWL[376] LDWL[375]
+ LDWL[374] LDWL[373] LDWL[372] LDWL[371] LDWL[370] LDWL[369] LDWL[368] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[3] LDL3X[5] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[22] LDWL[367] LDWL[366] LDWL[365] LDWL[364] LDWL[363] LDWL[362] LDWL[361] LDWL[360] LDWL[359]
+ LDWL[358] LDWL[357] LDWL[356] LDWL[355] LDWL[354] LDWL[353] LDWL[352] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[2] LDL3X[5] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[21] LDWL[351] LDWL[350] LDWL[349] LDWL[348] LDWL[347] LDWL[346] LDWL[345] LDWL[344] LDWL[343]
+ LDWL[342] LDWL[341] LDWL[340] LDWL[339] LDWL[338] LDWL[337] LDWL[336] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[1] LDL3X[5] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[20] LDWL[335] LDWL[334] LDWL[333] LDWL[332] LDWL[331] LDWL[330] LDWL[329] LDWL[328] LDWL[327]
+ LDWL[326] LDWL[325] LDWL[324] LDWL[323] LDWL[322] LDWL[321] LDWL[320] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[0] LDL3X[5] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[19] LDWL[319] LDWL[318] LDWL[317] LDWL[316] LDWL[315] LDWL[314] LDWL[313] LDWL[312] LDWL[311]
+ LDWL[310] LDWL[309] LDWL[308] LDWL[307] LDWL[306] LDWL[305] LDWL[304] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[3] LDL3X[4] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[18] LDWL[303] LDWL[302] LDWL[301] LDWL[300] LDWL[299] LDWL[298] LDWL[297] LDWL[296] LDWL[295]
+ LDWL[294] LDWL[293] LDWL[292] LDWL[291] LDWL[290] LDWL[289] LDWL[288] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[2] LDL3X[4] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[17] LDWL[287] LDWL[286] LDWL[285] LDWL[284] LDWL[283] LDWL[282] LDWL[281] LDWL[280] LDWL[279]
+ LDWL[278] LDWL[277] LDWL[276] LDWL[275] LDWL[274] LDWL[273] LDWL[272] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[1] LDL3X[4] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[16] LDWL[271] LDWL[270] LDWL[269] LDWL[268] LDWL[267] LDWL[266] LDWL[265] LDWL[264] LDWL[263]
+ LDWL[262] LDWL[261] LDWL[260] LDWL[259] LDWL[258] LDWL[257] LDWL[256] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[0] LDL3X[4] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[15] LDWL[255] LDWL[254] LDWL[253] LDWL[252] LDWL[251] LDWL[250] LDWL[249] LDWL[248] LDWL[247]
+ LDWL[246] LDWL[245] LDWL[244] LDWL[243] LDWL[242] LDWL[241] LDWL[240] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[3] LDL3X[3] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[14] LDWL[239] LDWL[238] LDWL[237] LDWL[236] LDWL[235] LDWL[234] LDWL[233] LDWL[232] LDWL[231]
+ LDWL[230] LDWL[229] LDWL[228] LDWL[227] LDWL[226] LDWL[225] LDWL[224] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[2] LDL3X[3] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[13] LDWL[223] LDWL[222] LDWL[221] LDWL[220] LDWL[219] LDWL[218] LDWL[217] LDWL[216] LDWL[215]
+ LDWL[214] LDWL[213] LDWL[212] LDWL[211] LDWL[210] LDWL[209] LDWL[208] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[1] LDL3X[3] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[12] LDWL[207] LDWL[206] LDWL[205] LDWL[204] LDWL[203] LDWL[202] LDWL[201] LDWL[200] LDWL[199]
+ LDWL[198] LDWL[197] LDWL[196] LDWL[195] LDWL[194] LDWL[193] LDWL[192] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[0] LDL3X[3] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[11] LDWL[191] LDWL[190] LDWL[189] LDWL[188] LDWL[187] LDWL[186] LDWL[185] LDWL[184] LDWL[183]
+ LDWL[182] LDWL[181] LDWL[180] LDWL[179] LDWL[178] LDWL[177] LDWL[176] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[3] LDL3X[2] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[10] LDWL[175] LDWL[174] LDWL[173] LDWL[172] LDWL[171] LDWL[170] LDWL[169] LDWL[168] LDWL[167]
+ LDWL[166] LDWL[165] LDWL[164] LDWL[163] LDWL[162] LDWL[161] LDWL[160] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[2] LDL3X[2] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[9] LDWL[159] LDWL[158] LDWL[157] LDWL[156] LDWL[155] LDWL[154] LDWL[153] LDWL[152] LDWL[151]
+ LDWL[150] LDWL[149] LDWL[148] LDWL[147] LDWL[146] LDWL[145] LDWL[144] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[1] LDL3X[2] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[8] LDWL[143] LDWL[142] LDWL[141] LDWL[140] LDWL[139] LDWL[138] LDWL[137] LDWL[136] LDWL[135]
+ LDWL[134] LDWL[133] LDWL[132] LDWL[131] LDWL[130] LDWL[129] LDWL[128] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[0] LDL3X[2] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[7] LDWL[127] LDWL[126] LDWL[125] LDWL[124] LDWL[123] LDWL[122] LDWL[121] LDWL[120] LDWL[119]
+ LDWL[118] LDWL[117] LDWL[116] LDWL[115] LDWL[114] LDWL[113] LDWL[112] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[3] LDL3X[1] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[6] LDWL[111] LDWL[110] LDWL[109] LDWL[108] LDWL[107] LDWL[106] LDWL[105] LDWL[104] LDWL[103]
+ LDWL[102] LDWL[101] LDWL[100] LDWL[99] LDWL[98] LDWL[97] LDWL[96] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12]
+ LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0]
+ LDL2X[2] LDL3X[1] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[5] LDWL[95] LDWL[94] LDWL[93] LDWL[92] LDWL[91] LDWL[90] LDWL[89] LDWL[88] LDWL[87] LDWL[86]
+ LDWL[85] LDWL[84] LDWL[83] LDWL[82] LDWL[81] LDWL[80] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12] LDL1X[11]
+ LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0] LDL2X[1]
+ LDL3X[1] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[4] LDWL[79] LDWL[78] LDWL[77] LDWL[76] LDWL[75] LDWL[74] LDWL[73] LDWL[72] LDWL[71] LDWL[70]
+ LDWL[69] LDWL[68] LDWL[67] LDWL[66] LDWL[65] LDWL[64] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12] LDL1X[11]
+ LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0] LDL2X[0]
+ LDL3X[1] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[3] LDWL[63] LDWL[62] LDWL[61] LDWL[60] LDWL[59] LDWL[58] LDWL[57] LDWL[56] LDWL[55] LDWL[54]
+ LDWL[53] LDWL[52] LDWL[51] LDWL[50] LDWL[49] LDWL[48] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12] LDL1X[11]
+ LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0] LDL2X[3]
+ LDL3X[0] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[2] LDWL[47] LDWL[46] LDWL[45] LDWL[44] LDWL[43] LDWL[42] LDWL[41] LDWL[40] LDWL[39] LDWL[38]
+ LDWL[37] LDWL[36] LDWL[35] LDWL[34] LDWL[33] LDWL[32] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12] LDL1X[11]
+ LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0] LDL2X[2]
+ LDL3X[0] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[1] LDWL[31] LDWL[30] LDWL[29] LDWL[28] LDWL[27] LDWL[26] LDWL[25] LDWL[24] LDWL[23] LDWL[22]
+ LDWL[21] LDWL[20] LDWL[19] LDWL[18] LDWL[17] LDWL[16] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12] LDL1X[11]
+ LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0] LDL2X[1]
+ LDL3X[0] LDCP_ROWDEC vss vccdec rom3_rowdec
xrdec[0] LDWL[15] LDWL[14] LDWL[13] LDWL[12] LDWL[11] LDWL[10] LDWL[9] LDWL[8] LDWL[7] LDWL[6]
+ LDWL[5] LDWL[4] LDWL[3] LDWL[2] LDWL[1] LDWL[0] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12] LDL1X[11] LDL1X[10]
+ LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0] LDL2X[0] LDL3X[0]
+ LDCP_ROWDEC vss vccdec rom3_rowdec
xrpre1 LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12] LDL1X[11] LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7]
+ LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0] LDAI[7] LDAI[6] LDAI[5] LDAI[4] vccdec vss
+ rom2_predec1
xrpre2 LDAI[12] LDAI[11] LDAI[10] LDAI[9] LDAI[8] vccdec vss LDL2X[3] LDL2X[2] LDL2X[1] LDL2X[0]
+ LDL3X[7] LDL3X[6] LDL3X[5] LDL3X[4] LDL3X[3] LDL3X[2] LDL3X[1] LDL3X[0] rom2_predec4
c3[7] LDL3X[7] vss 120f m=1
c3[6] LDL3X[6] vss 120f m=1
c3[5] LDL3X[5] vss 120f m=1
c3[4] LDL3X[4] vss 120f m=1
c3[3] LDL3X[3] vss 120f m=1
c3[2] LDL3X[2] vss 120f m=1
c3[1] LDL3X[1] vss 120f m=1
c3[0] LDL3X[0] vss 120f m=1
xcdecref LDYMSREF LDBLREF vccdec vss rom2_coldec_ref
xarr_ref LDWL[511] LDWL[510] LDWL[509] LDWL[508] LDWL[507] LDWL[506] LDWL[505] LDWL[504] LDWL[503]
+ LDWL[502] LDWL[501] LDWL[500] LDWL[499] LDWL[498] LDWL[497] LDWL[496] LDWL[495] LDWL[494] LDWL[493] LDWL[492]
+ LDWL[491] LDWL[490] LDWL[489] LDWL[488] LDWL[487] LDWL[486] LDWL[485] LDWL[484] LDWL[483] LDWL[482] LDWL[481]
+ LDWL[480] LDWL[479] LDWL[478] LDWL[477] LDWL[476] LDWL[475] LDWL[474] LDWL[473] LDWL[472] LDWL[471] LDWL[470]
+ LDWL[469] LDWL[468] LDWL[467] LDWL[466] LDWL[465] LDWL[464] LDWL[463] LDWL[462] LDWL[461] LDWL[460] LDWL[459]
+ LDWL[458] LDWL[457] LDWL[456] LDWL[455] LDWL[454] LDWL[453] LDWL[452] LDWL[451] LDWL[450] LDWL[449] LDWL[448]
+ LDWL[447] LDWL[446] LDWL[445] LDWL[444] LDWL[443] LDWL[442] LDWL[441] LDWL[440] LDWL[439] LDWL[438] LDWL[437]
+ LDWL[436] LDWL[435] LDWL[434] LDWL[433] LDWL[432] LDWL[431] LDWL[430] LDWL[429] LDWL[428] LDWL[427] LDWL[426]
+ LDWL[425] LDWL[424] LDWL[423] LDWL[422] LDWL[421] LDWL[420] LDWL[419] LDWL[418] LDWL[417] LDWL[416] LDWL[415]
+ LDWL[414] LDWL[413] LDWL[412] LDWL[411] LDWL[410] LDWL[409] LDWL[408] LDWL[407] LDWL[406] LDWL[405] LDWL[404]
+ LDWL[403] LDWL[402] LDWL[401] LDWL[400] LDWL[399] LDWL[398] LDWL[397] LDWL[396] LDWL[395] LDWL[394] LDWL[393]
+ LDWL[392] LDWL[391] LDWL[390] LDWL[389] LDWL[388] LDWL[387] LDWL[386] LDWL[385] LDWL[384] LDWL[383] LDWL[382]
+ LDWL[381] LDWL[380] LDWL[379] LDWL[378] LDWL[377] LDWL[376] LDWL[375] LDWL[374] LDWL[373] LDWL[372] LDWL[371]
+ LDWL[370] LDWL[369] LDWL[368] LDWL[367] LDWL[366] LDWL[365] LDWL[364] LDWL[363] LDWL[362] LDWL[361] LDWL[360]
+ LDWL[359] LDWL[358] LDWL[357] LDWL[356] LDWL[355] LDWL[354] LDWL[353] LDWL[352] LDWL[351] LDWL[350] LDWL[349]
+ LDWL[348] LDWL[347] LDWL[346] LDWL[345] LDWL[344] LDWL[343] LDWL[342] LDWL[341] LDWL[340] LDWL[339] LDWL[338]
+ LDWL[337] LDWL[336] LDWL[335] LDWL[334] LDWL[333] LDWL[332] LDWL[331] LDWL[330] LDWL[329] LDWL[328] LDWL[327]
+ LDWL[326] LDWL[325] LDWL[324] LDWL[323] LDWL[322] LDWL[321] LDWL[320] LDWL[319] LDWL[318] LDWL[317] LDWL[316]
+ LDWL[315] LDWL[314] LDWL[313] LDWL[312] LDWL[311] LDWL[310] LDWL[309] LDWL[308] LDWL[307] LDWL[306] LDWL[305]
+ LDWL[304] LDWL[303] LDWL[302] LDWL[301] LDWL[300] LDWL[299] LDWL[298] LDWL[297] LDWL[296] LDWL[295] LDWL[294]
+ LDWL[293] LDWL[292] LDWL[291] LDWL[290] LDWL[289] LDWL[288] LDWL[287] LDWL[286] LDWL[285] LDWL[284] LDWL[283]
+ LDWL[282] LDWL[281] LDWL[280] LDWL[279] LDWL[278] LDWL[277] LDWL[276] LDWL[275] LDWL[274] LDWL[273] LDWL[272]
+ LDWL[271] LDWL[270] LDWL[269] LDWL[268] LDWL[267] LDWL[266] LDWL[265] LDWL[264] LDWL[263] LDWL[262] LDWL[261]
+ LDWL[260] LDWL[259] LDWL[258] LDWL[257] LDWL[256] LDWL[255] LDWL[254] LDWL[253] LDWL[252] LDWL[251] LDWL[250]
+ LDWL[249] LDWL[248] LDWL[247] LDWL[246] LDWL[245] LDWL[244] LDWL[243] LDWL[242] LDWL[241] LDWL[240] LDWL[239]
+ LDWL[238] LDWL[237] LDWL[236] LDWL[235] LDWL[234] LDWL[233] LDWL[232] LDWL[231] LDWL[230] LDWL[229] LDWL[228]
+ LDWL[227] LDWL[226] LDWL[225] LDWL[224] LDWL[223] LDWL[222] LDWL[221] LDWL[220] LDWL[219] LDWL[218] LDWL[217]
+ LDWL[216] LDWL[215] LDWL[214] LDWL[213] LDWL[212] LDWL[211] LDWL[210] LDWL[209] LDWL[208] LDWL[207] LDWL[206]
+ LDWL[205] LDWL[204] LDWL[203] LDWL[202] LDWL[201] LDWL[200] LDWL[199] LDWL[198] LDWL[197] LDWL[196] LDWL[195]
+ LDWL[194] LDWL[193] LDWL[192] LDWL[191] LDWL[190] LDWL[189] LDWL[188] LDWL[187] LDWL[186] LDWL[185] LDWL[184]
+ LDWL[183] LDWL[182] LDWL[181] LDWL[180] LDWL[179] LDWL[178] LDWL[177] LDWL[176] LDWL[175] LDWL[174] LDWL[173]
+ LDWL[172] LDWL[171] LDWL[170] LDWL[169] LDWL[168] LDWL[167] LDWL[166] LDWL[165] LDWL[164] LDWL[163] LDWL[162]
+ LDWL[161] LDWL[160] LDWL[159] LDWL[158] LDWL[157] LDWL[156] LDWL[155] LDWL[154] LDWL[153] LDWL[152] LDWL[151]
+ LDWL[150] LDWL[149] LDWL[148] LDWL[147] LDWL[146] LDWL[145] LDWL[144] LDWL[143] LDWL[142] LDWL[141] LDWL[140]
+ LDWL[139] LDWL[138] LDWL[137] LDWL[136] LDWL[135] LDWL[134] LDWL[133] LDWL[132] LDWL[131] LDWL[130] LDWL[129]
+ LDWL[128] LDWL[127] LDWL[126] LDWL[125] LDWL[124] LDWL[123] LDWL[122] LDWL[121] LDWL[120] LDWL[119] LDWL[118]
+ LDWL[117] LDWL[116] LDWL[115] LDWL[114] LDWL[113] LDWL[112] LDWL[111] LDWL[110] LDWL[109] LDWL[108] LDWL[107]
+ LDWL[106] LDWL[105] LDWL[104] LDWL[103] LDWL[102] LDWL[101] LDWL[100] LDWL[99] LDWL[98] LDWL[97] LDWL[96]
+ LDWL[95] LDWL[94] LDWL[93] LDWL[92] LDWL[91] LDWL[90] LDWL[89] LDWL[88] LDWL[87] LDWL[86] LDWL[85] LDWL[84]
+ LDWL[83] LDWL[82] LDWL[81] LDWL[80] LDWL[79] LDWL[78] LDWL[77] LDWL[76] LDWL[75] LDWL[74] LDWL[73] LDWL[72]
+ LDWL[71] LDWL[70] LDWL[69] LDWL[68] LDWL[67] LDWL[66] LDWL[65] LDWL[64] LDWL[63] LDWL[62] LDWL[61] LDWL[60]
+ LDWL[59] LDWL[58] LDWL[57] LDWL[56] LDWL[55] LDWL[54] LDWL[53] LDWL[52] LDWL[51] LDWL[50] LDWL[49] LDWL[48]
+ LDWL[47] LDWL[46] LDWL[45] LDWL[44] LDWL[43] LDWL[42] LDWL[41] LDWL[40] LDWL[39] LDWL[38] LDWL[37] LDWL[36]
+ LDWL[35] LDWL[34] LDWL[33] LDWL[32] LDWL[31] LDWL[30] LDWL[29] LDWL[28] LDWL[27] LDWL[26] LDWL[25] LDWL[24]
+ LDWL[23] LDWL[22] LDWL[21] LDWL[20] LDWL[19] LDWL[18] LDWL[17] LDWL[16] LDWL[15] LDWL[14] LDWL[13] LDWL[12]
+ LDWL[11] LDWL[10] LDWL[9] LDWL[8] LDWL[7] LDWL[6] LDWL[5] LDWL[4] LDWL[3] LDWL[2] LDWL[1] LDWL[0] vss
+ LDBLREF rom3_array_ref
xcpr[256] LDCP_COL_B LDBL[255] vss rom2_col_prech
xcpr[255] LDCP_COL_B LDBL[254] vss rom2_col_prech
xcpr[254] LDCP_COL_B LDBL[253] vss rom2_col_prech
xcpr[253] LDCP_COL_B LDBL[252] vss rom2_col_prech
xcpr[252] LDCP_COL_B LDBL[251] vss rom2_col_prech
xcpr[251] LDCP_COL_B LDBL[250] vss rom2_col_prech
xcpr[250] LDCP_COL_B LDBL[249] vss rom2_col_prech
xcpr[249] LDCP_COL_B LDBL[248] vss rom2_col_prech
xcpr[248] LDCP_COL_B LDBL[247] vss rom2_col_prech
xcpr[247] LDCP_COL_B LDBL[246] vss rom2_col_prech
xcpr[246] LDCP_COL_B LDBL[245] vss rom2_col_prech
xcpr[245] LDCP_COL_B LDBL[244] vss rom2_col_prech
xcpr[244] LDCP_COL_B LDBL[243] vss rom2_col_prech
xcpr[243] LDCP_COL_B LDBL[242] vss rom2_col_prech
xcpr[242] LDCP_COL_B LDBL[241] vss rom2_col_prech
xcpr[241] LDCP_COL_B LDBL[240] vss rom2_col_prech
xcpr[240] LDCP_COL_B LDBL[239] vss rom2_col_prech
xcpr[239] LDCP_COL_B LDBL[238] vss rom2_col_prech
xcpr[238] LDCP_COL_B LDBL[237] vss rom2_col_prech
xcpr[237] LDCP_COL_B LDBL[236] vss rom2_col_prech
xcpr[236] LDCP_COL_B LDBL[235] vss rom2_col_prech
xcpr[235] LDCP_COL_B LDBL[234] vss rom2_col_prech
xcpr[234] LDCP_COL_B LDBL[233] vss rom2_col_prech
xcpr[233] LDCP_COL_B LDBL[232] vss rom2_col_prech
xcpr[232] LDCP_COL_B LDBL[231] vss rom2_col_prech
xcpr[231] LDCP_COL_B LDBL[230] vss rom2_col_prech
xcpr[230] LDCP_COL_B LDBL[229] vss rom2_col_prech
xcpr[229] LDCP_COL_B LDBL[228] vss rom2_col_prech
xcpr[228] LDCP_COL_B LDBL[227] vss rom2_col_prech
xcpr[227] LDCP_COL_B LDBL[226] vss rom2_col_prech
xcpr[226] LDCP_COL_B LDBL[225] vss rom2_col_prech
xcpr[225] LDCP_COL_B LDBL[224] vss rom2_col_prech
xcpr[224] LDCP_COL_B LDBL[223] vss rom2_col_prech
xcpr[223] LDCP_COL_B LDBL[222] vss rom2_col_prech
xcpr[222] LDCP_COL_B LDBL[221] vss rom2_col_prech
xcpr[221] LDCP_COL_B LDBL[220] vss rom2_col_prech
xcpr[220] LDCP_COL_B LDBL[219] vss rom2_col_prech
xcpr[219] LDCP_COL_B LDBL[218] vss rom2_col_prech
xcpr[218] LDCP_COL_B LDBL[217] vss rom2_col_prech
xcpr[217] LDCP_COL_B LDBL[216] vss rom2_col_prech
xcpr[216] LDCP_COL_B LDBL[215] vss rom2_col_prech
xcpr[215] LDCP_COL_B LDBL[214] vss rom2_col_prech
xcpr[214] LDCP_COL_B LDBL[213] vss rom2_col_prech
xcpr[213] LDCP_COL_B LDBL[212] vss rom2_col_prech
xcpr[212] LDCP_COL_B LDBL[211] vss rom2_col_prech
xcpr[211] LDCP_COL_B LDBL[210] vss rom2_col_prech
xcpr[210] LDCP_COL_B LDBL[209] vss rom2_col_prech
xcpr[209] LDCP_COL_B LDBL[208] vss rom2_col_prech
xcpr[208] LDCP_COL_B LDBL[207] vss rom2_col_prech
xcpr[207] LDCP_COL_B LDBL[206] vss rom2_col_prech
xcpr[206] LDCP_COL_B LDBL[205] vss rom2_col_prech
xcpr[205] LDCP_COL_B LDBL[204] vss rom2_col_prech
xcpr[204] LDCP_COL_B LDBL[203] vss rom2_col_prech
xcpr[203] LDCP_COL_B LDBL[202] vss rom2_col_prech
xcpr[202] LDCP_COL_B LDBL[201] vss rom2_col_prech
xcpr[201] LDCP_COL_B LDBL[200] vss rom2_col_prech
xcpr[200] LDCP_COL_B LDBL[199] vss rom2_col_prech
xcpr[199] LDCP_COL_B LDBL[198] vss rom2_col_prech
xcpr[198] LDCP_COL_B LDBL[197] vss rom2_col_prech
xcpr[197] LDCP_COL_B LDBL[196] vss rom2_col_prech
xcpr[196] LDCP_COL_B LDBL[195] vss rom2_col_prech
xcpr[195] LDCP_COL_B LDBL[194] vss rom2_col_prech
xcpr[194] LDCP_COL_B LDBL[193] vss rom2_col_prech
xcpr[193] LDCP_COL_B LDBL[192] vss rom2_col_prech
xcpr[192] LDCP_COL_B LDBL[191] vss rom2_col_prech
xcpr[191] LDCP_COL_B LDBL[190] vss rom2_col_prech
xcpr[190] LDCP_COL_B LDBL[189] vss rom2_col_prech
xcpr[189] LDCP_COL_B LDBL[188] vss rom2_col_prech
xcpr[188] LDCP_COL_B LDBL[187] vss rom2_col_prech
xcpr[187] LDCP_COL_B LDBL[186] vss rom2_col_prech
xcpr[186] LDCP_COL_B LDBL[185] vss rom2_col_prech
xcpr[185] LDCP_COL_B LDBL[184] vss rom2_col_prech
xcpr[184] LDCP_COL_B LDBL[183] vss rom2_col_prech
xcpr[183] LDCP_COL_B LDBL[182] vss rom2_col_prech
xcpr[182] LDCP_COL_B LDBL[181] vss rom2_col_prech
xcpr[181] LDCP_COL_B LDBL[180] vss rom2_col_prech
xcpr[180] LDCP_COL_B LDBL[179] vss rom2_col_prech
xcpr[179] LDCP_COL_B LDBL[178] vss rom2_col_prech
xcpr[178] LDCP_COL_B LDBL[177] vss rom2_col_prech
xcpr[177] LDCP_COL_B LDBL[176] vss rom2_col_prech
xcpr[176] LDCP_COL_B LDBL[175] vss rom2_col_prech
xcpr[175] LDCP_COL_B LDBL[174] vss rom2_col_prech
xcpr[174] LDCP_COL_B LDBL[173] vss rom2_col_prech
xcpr[173] LDCP_COL_B LDBL[172] vss rom2_col_prech
xcpr[172] LDCP_COL_B LDBL[171] vss rom2_col_prech
xcpr[171] LDCP_COL_B LDBL[170] vss rom2_col_prech
xcpr[170] LDCP_COL_B LDBL[169] vss rom2_col_prech
xcpr[169] LDCP_COL_B LDBL[168] vss rom2_col_prech
xcpr[168] LDCP_COL_B LDBL[167] vss rom2_col_prech
xcpr[167] LDCP_COL_B LDBL[166] vss rom2_col_prech
xcpr[166] LDCP_COL_B LDBL[165] vss rom2_col_prech
xcpr[165] LDCP_COL_B LDBL[164] vss rom2_col_prech
xcpr[164] LDCP_COL_B LDBL[163] vss rom2_col_prech
xcpr[163] LDCP_COL_B LDBL[162] vss rom2_col_prech
xcpr[162] LDCP_COL_B LDBL[161] vss rom2_col_prech
xcpr[161] LDCP_COL_B LDBL[160] vss rom2_col_prech
xcpr[160] LDCP_COL_B LDBL[159] vss rom2_col_prech
xcpr[159] LDCP_COL_B LDBL[158] vss rom2_col_prech
xcpr[158] LDCP_COL_B LDBL[157] vss rom2_col_prech
xcpr[157] LDCP_COL_B LDBL[156] vss rom2_col_prech
xcpr[156] LDCP_COL_B LDBL[155] vss rom2_col_prech
xcpr[155] LDCP_COL_B LDBL[154] vss rom2_col_prech
xcpr[154] LDCP_COL_B LDBL[153] vss rom2_col_prech
xcpr[153] LDCP_COL_B LDBL[152] vss rom2_col_prech
xcpr[152] LDCP_COL_B LDBL[151] vss rom2_col_prech
xcpr[151] LDCP_COL_B LDBL[150] vss rom2_col_prech
xcpr[150] LDCP_COL_B LDBL[149] vss rom2_col_prech
xcpr[149] LDCP_COL_B LDBL[148] vss rom2_col_prech
xcpr[148] LDCP_COL_B LDBL[147] vss rom2_col_prech
xcpr[147] LDCP_COL_B LDBL[146] vss rom2_col_prech
xcpr[146] LDCP_COL_B LDBL[145] vss rom2_col_prech
xcpr[145] LDCP_COL_B LDBL[144] vss rom2_col_prech
xcpr[144] LDCP_COL_B LDBL[143] vss rom2_col_prech
xcpr[143] LDCP_COL_B LDBL[142] vss rom2_col_prech
xcpr[142] LDCP_COL_B LDBL[141] vss rom2_col_prech
xcpr[141] LDCP_COL_B LDBL[140] vss rom2_col_prech
xcpr[140] LDCP_COL_B LDBL[139] vss rom2_col_prech
xcpr[139] LDCP_COL_B LDBL[138] vss rom2_col_prech
xcpr[138] LDCP_COL_B LDBL[137] vss rom2_col_prech
xcpr[137] LDCP_COL_B LDBL[136] vss rom2_col_prech
xcpr[136] LDCP_COL_B LDBL[135] vss rom2_col_prech
xcpr[135] LDCP_COL_B LDBL[134] vss rom2_col_prech
xcpr[134] LDCP_COL_B LDBL[133] vss rom2_col_prech
xcpr[133] LDCP_COL_B LDBL[132] vss rom2_col_prech
xcpr[132] LDCP_COL_B LDBL[131] vss rom2_col_prech
xcpr[131] LDCP_COL_B LDBL[130] vss rom2_col_prech
xcpr[130] LDCP_COL_B LDBL[129] vss rom2_col_prech
xcpr[129] LDCP_COL_B LDBL[128] vss rom2_col_prech
xcpr[128] LDCP_COL_B LDBL[127] vss rom2_col_prech
xcpr[127] LDCP_COL_B LDBL[126] vss rom2_col_prech
xcpr[126] LDCP_COL_B LDBL[125] vss rom2_col_prech
xcpr[125] LDCP_COL_B LDBL[124] vss rom2_col_prech
xcpr[124] LDCP_COL_B LDBL[123] vss rom2_col_prech
xcpr[123] LDCP_COL_B LDBL[122] vss rom2_col_prech
xcpr[122] LDCP_COL_B LDBL[121] vss rom2_col_prech
xcpr[121] LDCP_COL_B LDBL[120] vss rom2_col_prech
xcpr[120] LDCP_COL_B LDBL[119] vss rom2_col_prech
xcpr[119] LDCP_COL_B LDBL[118] vss rom2_col_prech
xcpr[118] LDCP_COL_B LDBL[117] vss rom2_col_prech
xcpr[117] LDCP_COL_B LDBL[116] vss rom2_col_prech
xcpr[116] LDCP_COL_B LDBL[115] vss rom2_col_prech
xcpr[115] LDCP_COL_B LDBL[114] vss rom2_col_prech
xcpr[114] LDCP_COL_B LDBL[113] vss rom2_col_prech
xcpr[113] LDCP_COL_B LDBL[112] vss rom2_col_prech
xcpr[112] LDCP_COL_B LDBL[111] vss rom2_col_prech
xcpr[111] LDCP_COL_B LDBL[110] vss rom2_col_prech
xcpr[110] LDCP_COL_B LDBL[109] vss rom2_col_prech
xcpr[109] LDCP_COL_B LDBL[108] vss rom2_col_prech
xcpr[108] LDCP_COL_B LDBL[107] vss rom2_col_prech
xcpr[107] LDCP_COL_B LDBL[106] vss rom2_col_prech
xcpr[106] LDCP_COL_B LDBL[105] vss rom2_col_prech
xcpr[105] LDCP_COL_B LDBL[104] vss rom2_col_prech
xcpr[104] LDCP_COL_B LDBL[103] vss rom2_col_prech
xcpr[103] LDCP_COL_B LDBL[102] vss rom2_col_prech
xcpr[102] LDCP_COL_B LDBL[101] vss rom2_col_prech
xcpr[101] LDCP_COL_B LDBL[100] vss rom2_col_prech
xcpr[100] LDCP_COL_B LDBL[99] vss rom2_col_prech
xcpr[99] LDCP_COL_B LDBL[98] vss rom2_col_prech
xcpr[98] LDCP_COL_B LDBL[97] vss rom2_col_prech
xcpr[97] LDCP_COL_B LDBL[96] vss rom2_col_prech
xcpr[96] LDCP_COL_B LDBL[95] vss rom2_col_prech
xcpr[95] LDCP_COL_B LDBL[94] vss rom2_col_prech
xcpr[94] LDCP_COL_B LDBL[93] vss rom2_col_prech
xcpr[93] LDCP_COL_B LDBL[92] vss rom2_col_prech
xcpr[92] LDCP_COL_B LDBL[91] vss rom2_col_prech
xcpr[91] LDCP_COL_B LDBL[90] vss rom2_col_prech
xcpr[90] LDCP_COL_B LDBL[89] vss rom2_col_prech
xcpr[89] LDCP_COL_B LDBL[88] vss rom2_col_prech
xcpr[88] LDCP_COL_B LDBL[87] vss rom2_col_prech
xcpr[87] LDCP_COL_B LDBL[86] vss rom2_col_prech
xcpr[86] LDCP_COL_B LDBL[85] vss rom2_col_prech
xcpr[85] LDCP_COL_B LDBL[84] vss rom2_col_prech
xcpr[84] LDCP_COL_B LDBL[83] vss rom2_col_prech
xcpr[83] LDCP_COL_B LDBL[82] vss rom2_col_prech
xcpr[82] LDCP_COL_B LDBL[81] vss rom2_col_prech
xcpr[81] LDCP_COL_B LDBL[80] vss rom2_col_prech
xcpr[80] LDCP_COL_B LDBL[79] vss rom2_col_prech
xcpr[79] LDCP_COL_B LDBL[78] vss rom2_col_prech
xcpr[78] LDCP_COL_B LDBL[77] vss rom2_col_prech
xcpr[77] LDCP_COL_B LDBL[76] vss rom2_col_prech
xcpr[76] LDCP_COL_B LDBL[75] vss rom2_col_prech
xcpr[75] LDCP_COL_B LDBL[74] vss rom2_col_prech
xcpr[74] LDCP_COL_B LDBL[73] vss rom2_col_prech
xcpr[73] LDCP_COL_B LDBL[72] vss rom2_col_prech
xcpr[72] LDCP_COL_B LDBL[71] vss rom2_col_prech
xcpr[71] LDCP_COL_B LDBL[70] vss rom2_col_prech
xcpr[70] LDCP_COL_B LDBL[69] vss rom2_col_prech
xcpr[69] LDCP_COL_B LDBL[68] vss rom2_col_prech
xcpr[68] LDCP_COL_B LDBL[67] vss rom2_col_prech
xcpr[67] LDCP_COL_B LDBL[66] vss rom2_col_prech
xcpr[66] LDCP_COL_B LDBL[65] vss rom2_col_prech
xcpr[65] LDCP_COL_B LDBL[64] vss rom2_col_prech
xcpr[64] LDCP_COL_B LDBL[63] vss rom2_col_prech
xcpr[63] LDCP_COL_B LDBL[62] vss rom2_col_prech
xcpr[62] LDCP_COL_B LDBL[61] vss rom2_col_prech
xcpr[61] LDCP_COL_B LDBL[60] vss rom2_col_prech
xcpr[60] LDCP_COL_B LDBL[59] vss rom2_col_prech
xcpr[59] LDCP_COL_B LDBL[58] vss rom2_col_prech
xcpr[58] LDCP_COL_B LDBL[57] vss rom2_col_prech
xcpr[57] LDCP_COL_B LDBL[56] vss rom2_col_prech
xcpr[56] LDCP_COL_B LDBL[55] vss rom2_col_prech
xcpr[55] LDCP_COL_B LDBL[54] vss rom2_col_prech
xcpr[54] LDCP_COL_B LDBL[53] vss rom2_col_prech
xcpr[53] LDCP_COL_B LDBL[52] vss rom2_col_prech
xcpr[52] LDCP_COL_B LDBL[51] vss rom2_col_prech
xcpr[51] LDCP_COL_B LDBL[50] vss rom2_col_prech
xcpr[50] LDCP_COL_B LDBL[49] vss rom2_col_prech
xcpr[49] LDCP_COL_B LDBL[48] vss rom2_col_prech
xcpr[48] LDCP_COL_B LDBL[47] vss rom2_col_prech
xcpr[47] LDCP_COL_B LDBL[46] vss rom2_col_prech
xcpr[46] LDCP_COL_B LDBL[45] vss rom2_col_prech
xcpr[45] LDCP_COL_B LDBL[44] vss rom2_col_prech
xcpr[44] LDCP_COL_B LDBL[43] vss rom2_col_prech
xcpr[43] LDCP_COL_B LDBL[42] vss rom2_col_prech
xcpr[42] LDCP_COL_B LDBL[41] vss rom2_col_prech
xcpr[41] LDCP_COL_B LDBL[40] vss rom2_col_prech
xcpr[40] LDCP_COL_B LDBL[39] vss rom2_col_prech
xcpr[39] LDCP_COL_B LDBL[38] vss rom2_col_prech
xcpr[38] LDCP_COL_B LDBL[37] vss rom2_col_prech
xcpr[37] LDCP_COL_B LDBL[36] vss rom2_col_prech
xcpr[36] LDCP_COL_B LDBL[35] vss rom2_col_prech
xcpr[35] LDCP_COL_B LDBL[34] vss rom2_col_prech
xcpr[34] LDCP_COL_B LDBL[33] vss rom2_col_prech
xcpr[33] LDCP_COL_B LDBL[32] vss rom2_col_prech
xcpr[32] LDCP_COL_B LDBL[31] vss rom2_col_prech
xcpr[31] LDCP_COL_B LDBL[30] vss rom2_col_prech
xcpr[30] LDCP_COL_B LDBL[29] vss rom2_col_prech
xcpr[29] LDCP_COL_B LDBL[28] vss rom2_col_prech
xcpr[28] LDCP_COL_B LDBL[27] vss rom2_col_prech
xcpr[27] LDCP_COL_B LDBL[26] vss rom2_col_prech
xcpr[26] LDCP_COL_B LDBL[25] vss rom2_col_prech
xcpr[25] LDCP_COL_B LDBL[24] vss rom2_col_prech
xcpr[24] LDCP_COL_B LDBL[23] vss rom2_col_prech
xcpr[23] LDCP_COL_B LDBL[22] vss rom2_col_prech
xcpr[22] LDCP_COL_B LDBL[21] vss rom2_col_prech
xcpr[21] LDCP_COL_B LDBL[20] vss rom2_col_prech
xcpr[20] LDCP_COL_B LDBL[19] vss rom2_col_prech
xcpr[19] LDCP_COL_B LDBL[18] vss rom2_col_prech
xcpr[18] LDCP_COL_B LDBL[17] vss rom2_col_prech
xcpr[17] LDCP_COL_B LDBL[16] vss rom2_col_prech
xcpr[16] LDCP_COL_B LDBL[15] vss rom2_col_prech
xcpr[15] LDCP_COL_B LDBL[14] vss rom2_col_prech
xcpr[14] LDCP_COL_B LDBL[13] vss rom2_col_prech
xcpr[13] LDCP_COL_B LDBL[12] vss rom2_col_prech
xcpr[12] LDCP_COL_B LDBL[11] vss rom2_col_prech
xcpr[11] LDCP_COL_B LDBL[10] vss rom2_col_prech
xcpr[10] LDCP_COL_B LDBL[9] vss rom2_col_prech
xcpr[9] LDCP_COL_B LDBL[8] vss rom2_col_prech
xcpr[8] LDCP_COL_B LDBL[7] vss rom2_col_prech
xcpr[7] LDCP_COL_B LDBL[6] vss rom2_col_prech
xcpr[6] LDCP_COL_B LDBL[5] vss rom2_col_prech
xcpr[5] LDCP_COL_B LDBL[4] vss rom2_col_prech
xcpr[4] LDCP_COL_B LDBL[3] vss rom2_col_prech
xcpr[3] LDCP_COL_B LDBL[2] vss rom2_col_prech
xcpr[2] LDCP_COL_B LDBL[1] vss rom2_col_prech
xcpr[1] LDCP_COL_B LDBL[0] vss rom2_col_prech
xcpr[0] LDCP_COL_B LDBLREF vss rom2_col_prech
c0 LDPRECH vss 66f m=1
c6 LDSAL vss 34f m=1
c7 LDCP_ROWDEC vss 280f m=1
c8 LDCP_SA vss 44f m=1
c9 LDCP_COL_B vss 63f m=1
c10 LDCP_ADDLAT_B vss 12f m=1
.save  v(ldq[15])
.save  v(ldq[14])
.save  v(ldq[13])
.save  v(ldq[12])
.save  v(ldq[11])
.save  v(ldq[10])
.save  v(ldq[9])
.save  v(ldq[8])
.save  v(ldq[7])
.save  v(ldq[6])
.save  v(ldq[5])
.save  v(ldq[4])
.save  v(ldq[3])
.save  v(ldq[2])
.save  v(ldq[1])
.save  v(ldq[0])
.save  v(ldl1x[15])
.save  v(ldl1x[14])
.save  v(ldl1x[13])
.save  v(ldl1x[12])
.save  v(ldl1x[11])
.save  v(ldl1x[10])
.save  v(ldl1x[9])
.save  v(ldl1x[8])
.save  v(ldl1x[7])
.save  v(ldl1x[6])
.save  v(ldl1x[5])
.save  v(ldl1x[4])
.save  v(ldl1x[3])
.save  v(ldl1x[2])
.save  v(ldl1x[1])
.save  v(ldl1x[0])
.save  v(ldy1[15])
.save  v(ldy1[14])
.save  v(ldy1[13])
.save  v(ldy1[12])
.save  v(ldy1[11])
.save  v(ldy1[10])
.save  v(ldy1[9])
.save  v(ldy1[8])
.save  v(ldy1[7])
.save  v(ldy1[6])
.save  v(ldy1[5])
.save  v(ldy1[4])
.save  v(ldy1[3])
.save  v(ldy1[2])
.save  v(ldy1[1])
.save  v(ldy1[0])
.save  v(ldl3x[7])
.save  v(ldl3x[6])
.save  v(ldl3x[5])
.save  v(ldl3x[4])
.save  v(ldl3x[3])
.save  v(ldl3x[2])
.save  v(ldl3x[1])
.save  v(ldl3x[0])
.save  v(ldl2x[3])
.save  v(ldl2x[2])
.save  v(ldl2x[1])
.save  v(ldl2x[0])
.save  v(ldai[12])
.save  v(ldai[11])
.save  v(ldai[10])
.save  v(ldai[9])
.save  v(ldai[8])
.save  v(ldai[7])
.save  v(ldai[6])
.save  v(ldai[5])
.save  v(ldai[4])
.save  v(ldai[3])
.save  v(ldai[2])
.save  v(ldai[1])
.save  v(ldai[0])
.save  v(ldcp_sa)
.save  v(ldcp_rowdec)
.save  v(ldcp_addlat_b)
.save  v(ldcp_col_b)
.save  v(ldprech)
.save  v(ldsal)
.save  v(ldymsref)
.save  v(lden_lat)
.save  v(ldblref)
.save  v(ldyms[15])
.save  v(ldyms[14])
.save  v(ldyms[13])
.save  v(ldyms[12])
.save  v(ldyms[11])
.save  v(ldyms[10])
.save  v(ldyms[9])
.save  v(ldyms[8])
.save  v(ldyms[7])
.save  v(ldyms[6])
.save  v(ldyms[5])
.save  v(ldyms[4])
.save  v(ldyms[3])
.save  v(ldyms[2])
.save  v(ldyms[1])
.save  v(ldyms[0])
.save  v(ldoe)
.save  v(ldcp)
.save  v(lden)
.save  v(lda[12])
.save  v(lda[11])
.save  v(lda[10])
.save  v(lda[9])
.save  v(lda[8])
.save  v(lda[7])
.save  v(lda[6])
.save  v(lda[5])
.save  v(lda[4])
.save  v(lda[3])
.save  v(lda[2])
.save  v(lda[1])
.save  v(lda[0])
xarr LDWL[511] LDWL[510] LDWL[509] LDWL[508] LDWL[507] LDWL[506] LDWL[505] LDWL[504] LDWL[503]
+ LDWL[502] LDWL[501] LDWL[500] LDWL[499] LDWL[498] LDWL[497] LDWL[496] LDWL[495] LDWL[494] LDWL[493] LDWL[492]
+ LDWL[491] LDWL[490] LDWL[489] LDWL[488] LDWL[487] LDWL[486] LDWL[485] LDWL[484] LDWL[483] LDWL[482] LDWL[481]
+ LDWL[480] LDWL[479] LDWL[478] LDWL[477] LDWL[476] LDWL[475] LDWL[474] LDWL[473] LDWL[472] LDWL[471] LDWL[470]
+ LDWL[469] LDWL[468] LDWL[467] LDWL[466] LDWL[465] LDWL[464] LDWL[463] LDWL[462] LDWL[461] LDWL[460] LDWL[459]
+ LDWL[458] LDWL[457] LDWL[456] LDWL[455] LDWL[454] LDWL[453] LDWL[452] LDWL[451] LDWL[450] LDWL[449] LDWL[448]
+ LDWL[447] LDWL[446] LDWL[445] LDWL[444] LDWL[443] LDWL[442] LDWL[441] LDWL[440] LDWL[439] LDWL[438] LDWL[437]
+ LDWL[436] LDWL[435] LDWL[434] LDWL[433] LDWL[432] LDWL[431] LDWL[430] LDWL[429] LDWL[428] LDWL[427] LDWL[426]
+ LDWL[425] LDWL[424] LDWL[423] LDWL[422] LDWL[421] LDWL[420] LDWL[419] LDWL[418] LDWL[417] LDWL[416] LDWL[415]
+ LDWL[414] LDWL[413] LDWL[412] LDWL[411] LDWL[410] LDWL[409] LDWL[408] LDWL[407] LDWL[406] LDWL[405] LDWL[404]
+ LDWL[403] LDWL[402] LDWL[401] LDWL[400] LDWL[399] LDWL[398] LDWL[397] LDWL[396] LDWL[395] LDWL[394] LDWL[393]
+ LDWL[392] LDWL[391] LDWL[390] LDWL[389] LDWL[388] LDWL[387] LDWL[386] LDWL[385] LDWL[384] LDWL[383] LDWL[382]
+ LDWL[381] LDWL[380] LDWL[379] LDWL[378] LDWL[377] LDWL[376] LDWL[375] LDWL[374] LDWL[373] LDWL[372] LDWL[371]
+ LDWL[370] LDWL[369] LDWL[368] LDWL[367] LDWL[366] LDWL[365] LDWL[364] LDWL[363] LDWL[362] LDWL[361] LDWL[360]
+ LDWL[359] LDWL[358] LDWL[357] LDWL[356] LDWL[355] LDWL[354] LDWL[353] LDWL[352] LDWL[351] LDWL[350] LDWL[349]
+ LDWL[348] LDWL[347] LDWL[346] LDWL[345] LDWL[344] LDWL[343] LDWL[342] LDWL[341] LDWL[340] LDWL[339] LDWL[338]
+ LDWL[337] LDWL[336] LDWL[335] LDWL[334] LDWL[333] LDWL[332] LDWL[331] LDWL[330] LDWL[329] LDWL[328] LDWL[327]
+ LDWL[326] LDWL[325] LDWL[324] LDWL[323] LDWL[322] LDWL[321] LDWL[320] LDWL[319] LDWL[318] LDWL[317] LDWL[316]
+ LDWL[315] LDWL[314] LDWL[313] LDWL[312] LDWL[311] LDWL[310] LDWL[309] LDWL[308] LDWL[307] LDWL[306] LDWL[305]
+ LDWL[304] LDWL[303] LDWL[302] LDWL[301] LDWL[300] LDWL[299] LDWL[298] LDWL[297] LDWL[296] LDWL[295] LDWL[294]
+ LDWL[293] LDWL[292] LDWL[291] LDWL[290] LDWL[289] LDWL[288] LDWL[287] LDWL[286] LDWL[285] LDWL[284] LDWL[283]
+ LDWL[282] LDWL[281] LDWL[280] LDWL[279] LDWL[278] LDWL[277] LDWL[276] LDWL[275] LDWL[274] LDWL[273] LDWL[272]
+ LDWL[271] LDWL[270] LDWL[269] LDWL[268] LDWL[267] LDWL[266] LDWL[265] LDWL[264] LDWL[263] LDWL[262] LDWL[261]
+ LDWL[260] LDWL[259] LDWL[258] LDWL[257] LDWL[256] LDWL[255] LDWL[254] LDWL[253] LDWL[252] LDWL[251] LDWL[250]
+ LDWL[249] LDWL[248] LDWL[247] LDWL[246] LDWL[245] LDWL[244] LDWL[243] LDWL[242] LDWL[241] LDWL[240] LDWL[239]
+ LDWL[238] LDWL[237] LDWL[236] LDWL[235] LDWL[234] LDWL[233] LDWL[232] LDWL[231] LDWL[230] LDWL[229] LDWL[228]
+ LDWL[227] LDWL[226] LDWL[225] LDWL[224] LDWL[223] LDWL[222] LDWL[221] LDWL[220] LDWL[219] LDWL[218] LDWL[217]
+ LDWL[216] LDWL[215] LDWL[214] LDWL[213] LDWL[212] LDWL[211] LDWL[210] LDWL[209] LDWL[208] LDWL[207] LDWL[206]
+ LDWL[205] LDWL[204] LDWL[203] LDWL[202] LDWL[201] LDWL[200] LDWL[199] LDWL[198] LDWL[197] LDWL[196] LDWL[195]
+ LDWL[194] LDWL[193] LDWL[192] LDWL[191] LDWL[190] LDWL[189] LDWL[188] LDWL[187] LDWL[186] LDWL[185] LDWL[184]
+ LDWL[183] LDWL[182] LDWL[181] LDWL[180] LDWL[179] LDWL[178] LDWL[177] LDWL[176] LDWL[175] LDWL[174] LDWL[173]
+ LDWL[172] LDWL[171] LDWL[170] LDWL[169] LDWL[168] LDWL[167] LDWL[166] LDWL[165] LDWL[164] LDWL[163] LDWL[162]
+ LDWL[161] LDWL[160] LDWL[159] LDWL[158] LDWL[157] LDWL[156] LDWL[155] LDWL[154] LDWL[153] LDWL[152] LDWL[151]
+ LDWL[150] LDWL[149] LDWL[148] LDWL[147] LDWL[146] LDWL[145] LDWL[144] LDWL[143] LDWL[142] LDWL[141] LDWL[140]
+ LDWL[139] LDWL[138] LDWL[137] LDWL[136] LDWL[135] LDWL[134] LDWL[133] LDWL[132] LDWL[131] LDWL[130] LDWL[129]
+ LDWL[128] LDWL[127] LDWL[126] LDWL[125] LDWL[124] LDWL[123] LDWL[122] LDWL[121] LDWL[120] LDWL[119] LDWL[118]
+ LDWL[117] LDWL[116] LDWL[115] LDWL[114] LDWL[113] LDWL[112] LDWL[111] LDWL[110] LDWL[109] LDWL[108] LDWL[107]
+ LDWL[106] LDWL[105] LDWL[104] LDWL[103] LDWL[102] LDWL[101] LDWL[100] LDWL[99] LDWL[98] LDWL[97] LDWL[96]
+ LDWL[95] LDWL[94] LDWL[93] LDWL[92] LDWL[91] LDWL[90] LDWL[89] LDWL[88] LDWL[87] LDWL[86] LDWL[85] LDWL[84]
+ LDWL[83] LDWL[82] LDWL[81] LDWL[80] LDWL[79] LDWL[78] LDWL[77] LDWL[76] LDWL[75] LDWL[74] LDWL[73] LDWL[72]
+ LDWL[71] LDWL[70] LDWL[69] LDWL[68] LDWL[67] LDWL[66] LDWL[65] LDWL[64] LDWL[63] LDWL[62] LDWL[61] LDWL[60]
+ LDWL[59] LDWL[58] LDWL[57] LDWL[56] LDWL[55] LDWL[54] LDWL[53] LDWL[52] LDWL[51] LDWL[50] LDWL[49] LDWL[48]
+ LDWL[47] LDWL[46] LDWL[45] LDWL[44] LDWL[43] LDWL[42] LDWL[41] LDWL[40] LDWL[39] LDWL[38] LDWL[37] LDWL[36]
+ LDWL[35] LDWL[34] LDWL[33] LDWL[32] LDWL[31] LDWL[30] LDWL[29] LDWL[28] LDWL[27] LDWL[26] LDWL[25] LDWL[24]
+ LDWL[23] LDWL[22] LDWL[21] LDWL[20] LDWL[19] LDWL[18] LDWL[17] LDWL[16] LDWL[15] LDWL[14] LDWL[13] LDWL[12]
+ LDWL[11] LDWL[10] LDWL[9] LDWL[8] LDWL[7] LDWL[6] LDWL[5] LDWL[4] LDWL[3] LDWL[2] LDWL[1] LDWL[0] LDBL[255]
+ LDBL[254] LDBL[253] LDBL[252] LDBL[251] LDBL[250] LDBL[249] LDBL[248] LDBL[247] LDBL[246] LDBL[245] LDBL[244]
+ LDBL[243] LDBL[242] LDBL[241] LDBL[240] LDBL[239] LDBL[238] LDBL[237] LDBL[236] LDBL[235] LDBL[234] LDBL[233]
+ LDBL[232] LDBL[231] LDBL[230] LDBL[229] LDBL[228] LDBL[227] LDBL[226] LDBL[225] LDBL[224] LDBL[223] LDBL[222]
+ LDBL[221] LDBL[220] LDBL[219] LDBL[218] LDBL[217] LDBL[216] LDBL[215] LDBL[214] LDBL[213] LDBL[212] LDBL[211]
+ LDBL[210] LDBL[209] LDBL[208] LDBL[207] LDBL[206] LDBL[205] LDBL[204] LDBL[203] LDBL[202] LDBL[201] LDBL[200]
+ LDBL[199] LDBL[198] LDBL[197] LDBL[196] LDBL[195] LDBL[194] LDBL[193] LDBL[192] LDBL[191] LDBL[190] LDBL[189]
+ LDBL[188] LDBL[187] LDBL[186] LDBL[185] LDBL[184] LDBL[183] LDBL[182] LDBL[181] LDBL[180] LDBL[179] LDBL[178]
+ LDBL[177] LDBL[176] LDBL[175] LDBL[174] LDBL[173] LDBL[172] LDBL[171] LDBL[170] LDBL[169] LDBL[168] LDBL[167]
+ LDBL[166] LDBL[165] LDBL[164] LDBL[163] LDBL[162] LDBL[161] LDBL[160] LDBL[159] LDBL[158] LDBL[157] LDBL[156]
+ LDBL[155] LDBL[154] LDBL[153] LDBL[152] LDBL[151] LDBL[150] LDBL[149] LDBL[148] LDBL[147] LDBL[146] LDBL[145]
+ LDBL[144] LDBL[143] LDBL[142] LDBL[141] LDBL[140] LDBL[139] LDBL[138] LDBL[137] LDBL[136] LDBL[135] LDBL[134]
+ LDBL[133] LDBL[132] LDBL[131] LDBL[130] LDBL[129] LDBL[128] LDBL[127] LDBL[126] LDBL[125] LDBL[124] LDBL[123]
+ LDBL[122] LDBL[121] LDBL[120] LDBL[119] LDBL[118] LDBL[117] LDBL[116] LDBL[115] LDBL[114] LDBL[113] LDBL[112]
+ LDBL[111] LDBL[110] LDBL[109] LDBL[108] LDBL[107] LDBL[106] LDBL[105] LDBL[104] LDBL[103] LDBL[102] LDBL[101]
+ LDBL[100] LDBL[99] LDBL[98] LDBL[97] LDBL[96] LDBL[95] LDBL[94] LDBL[93] LDBL[92] LDBL[91] LDBL[90] LDBL[89]
+ LDBL[88] LDBL[87] LDBL[86] LDBL[85] LDBL[84] LDBL[83] LDBL[82] LDBL[81] LDBL[80] LDBL[79] LDBL[78] LDBL[77]
+ LDBL[76] LDBL[75] LDBL[74] LDBL[73] LDBL[72] LDBL[71] LDBL[70] LDBL[69] LDBL[68] LDBL[67] LDBL[66] LDBL[65]
+ LDBL[64] LDBL[63] LDBL[62] LDBL[61] LDBL[60] LDBL[59] LDBL[58] LDBL[57] LDBL[56] LDBL[55] LDBL[54] LDBL[53]
+ LDBL[52] LDBL[51] LDBL[50] LDBL[49] LDBL[48] LDBL[47] LDBL[46] LDBL[45] LDBL[44] LDBL[43] LDBL[42] LDBL[41]
+ LDBL[40] LDBL[39] LDBL[38] LDBL[37] LDBL[36] LDBL[35] LDBL[34] LDBL[33] LDBL[32] LDBL[31] LDBL[30] LDBL[29]
+ LDBL[28] LDBL[27] LDBL[26] LDBL[25] LDBL[24] LDBL[23] LDBL[22] LDBL[21] LDBL[20] LDBL[19] LDBL[18] LDBL[17]
+ LDBL[16] LDBL[15] LDBL[14] LDBL[13] LDBL[12] LDBL[11] LDBL[10] LDBL[9] LDBL[8] LDBL[7] LDBL[6] LDBL[5]
+ LDBL[4] LDBL[3] LDBL[2] LDBL[1] LDBL[0] vss rom3_array
.save  v(ldymsref)
.save  v(vcc)
.save  v(ldwl[511])
.save  v(ldwl[510])
.save  v(ldwl[509])
.save  v(ldwl[508])
.save  v(ldwl[507])
.save  v(ldwl[506])
.save  v(ldwl[505])
.save  v(ldwl[504])
.save  v(ldwl[503])
.save  v(ldwl[502])
.save  v(ldwl[501])
.save  v(ldwl[500])
.save  v(ldwl[499])
.save  v(ldwl[498])
.save  v(ldwl[497])
.save  v(ldwl[496])
.save  v(ldwl[495])
.save  v(ldwl[494])
.save  v(ldwl[493])
.save  v(ldwl[492])
.save  v(ldwl[491])
.save  v(ldwl[490])
.save  v(ldwl[489])
.save  v(ldwl[488])
.save  v(ldwl[487])
.save  v(ldwl[486])
.save  v(ldwl[485])
.save  v(ldwl[484])
.save  v(ldwl[483])
.save  v(ldwl[482])
.save  v(ldwl[481])
.save  v(ldwl[480])
.save  v(ldwl[479])
.save  v(ldwl[478])
.save  v(ldwl[477])
.save  v(ldwl[476])
.save  v(ldwl[475])
.save  v(ldwl[474])
.save  v(ldwl[473])
.save  v(ldwl[472])
.save  v(ldwl[471])
.save  v(ldwl[470])
.save  v(ldwl[469])
.save  v(ldwl[468])
.save  v(ldwl[467])
.save  v(ldwl[466])
.save  v(ldwl[465])
.save  v(ldwl[464])
.save  v(ldwl[463])
.save  v(ldwl[462])
.save  v(ldwl[461])
.save  v(ldwl[460])
.save  v(ldwl[459])
.save  v(ldwl[458])
.save  v(ldwl[457])
.save  v(ldwl[456])
.save  v(ldwl[455])
.save  v(ldwl[454])
.save  v(ldwl[453])
.save  v(ldwl[452])
.save  v(ldwl[451])
.save  v(ldwl[450])
.save  v(ldwl[449])
.save  v(ldwl[448])
.save  v(ldwl[447])
.save  v(ldwl[446])
.save  v(ldwl[445])
.save  v(ldwl[444])
.save  v(ldwl[443])
.save  v(ldwl[442])
.save  v(ldwl[441])
.save  v(ldwl[440])
.save  v(ldwl[439])
.save  v(ldwl[438])
.save  v(ldwl[437])
.save  v(ldwl[436])
.save  v(ldwl[435])
.save  v(ldwl[434])
.save  v(ldwl[433])
.save  v(ldwl[432])
.save  v(ldwl[431])
.save  v(ldwl[430])
.save  v(ldwl[429])
.save  v(ldwl[428])
.save  v(ldwl[427])
.save  v(ldwl[426])
.save  v(ldwl[425])
.save  v(ldwl[424])
.save  v(ldwl[423])
.save  v(ldwl[422])
.save  v(ldwl[421])
.save  v(ldwl[420])
.save  v(ldwl[419])
.save  v(ldwl[418])
.save  v(ldwl[417])
.save  v(ldwl[416])
.save  v(ldwl[415])
.save  v(ldwl[414])
.save  v(ldwl[413])
.save  v(ldwl[412])
.save  v(ldwl[411])
.save  v(ldwl[410])
.save  v(ldwl[409])
.save  v(ldwl[408])
.save  v(ldwl[407])
.save  v(ldwl[406])
.save  v(ldwl[405])
.save  v(ldwl[404])
.save  v(ldwl[403])
.save  v(ldwl[402])
.save  v(ldwl[401])
.save  v(ldwl[400])
.save  v(ldwl[399])
.save  v(ldwl[398])
.save  v(ldwl[397])
.save  v(ldwl[396])
.save  v(ldwl[395])
.save  v(ldwl[394])
.save  v(ldwl[393])
.save  v(ldwl[392])
.save  v(ldwl[391])
.save  v(ldwl[390])
.save  v(ldwl[389])
.save  v(ldwl[388])
.save  v(ldwl[387])
.save  v(ldwl[386])
.save  v(ldwl[385])
.save  v(ldwl[384])
.save  v(ldwl[383])
.save  v(ldwl[382])
.save  v(ldwl[381])
.save  v(ldwl[380])
.save  v(ldwl[379])
.save  v(ldwl[378])
.save  v(ldwl[377])
.save  v(ldwl[376])
.save  v(ldwl[375])
.save  v(ldwl[374])
.save  v(ldwl[373])
.save  v(ldwl[372])
.save  v(ldwl[371])
.save  v(ldwl[370])
.save  v(ldwl[369])
.save  v(ldwl[368])
.save  v(ldwl[367])
.save  v(ldwl[366])
.save  v(ldwl[365])
.save  v(ldwl[364])
.save  v(ldwl[363])
.save  v(ldwl[362])
.save  v(ldwl[361])
.save  v(ldwl[360])
.save  v(ldwl[359])
.save  v(ldwl[358])
.save  v(ldwl[357])
.save  v(ldwl[356])
.save  v(ldwl[355])
.save  v(ldwl[354])
.save  v(ldwl[353])
.save  v(ldwl[352])
.save  v(ldwl[351])
.save  v(ldwl[350])
.save  v(ldwl[349])
.save  v(ldwl[348])
.save  v(ldwl[347])
.save  v(ldwl[346])
.save  v(ldwl[345])
.save  v(ldwl[344])
.save  v(ldwl[343])
.save  v(ldwl[342])
.save  v(ldwl[341])
.save  v(ldwl[340])
.save  v(ldwl[339])
.save  v(ldwl[338])
.save  v(ldwl[337])
.save  v(ldwl[336])
.save  v(ldwl[335])
.save  v(ldwl[334])
.save  v(ldwl[333])
.save  v(ldwl[332])
.save  v(ldwl[331])
.save  v(ldwl[330])
.save  v(ldwl[329])
.save  v(ldwl[328])
.save  v(ldwl[327])
.save  v(ldwl[326])
.save  v(ldwl[325])
.save  v(ldwl[324])
.save  v(ldwl[323])
.save  v(ldwl[322])
.save  v(ldwl[321])
.save  v(ldwl[320])
.save  v(ldwl[319])
.save  v(ldwl[318])
.save  v(ldwl[317])
.save  v(ldwl[316])
.save  v(ldwl[315])
.save  v(ldwl[314])
.save  v(ldwl[313])
.save  v(ldwl[312])
.save  v(ldwl[311])
.save  v(ldwl[310])
.save  v(ldwl[309])
.save  v(ldwl[308])
.save  v(ldwl[307])
.save  v(ldwl[306])
.save  v(ldwl[305])
.save  v(ldwl[304])
.save  v(ldwl[303])
.save  v(ldwl[302])
.save  v(ldwl[301])
.save  v(ldwl[300])
.save  v(ldwl[299])
.save  v(ldwl[298])
.save  v(ldwl[297])
.save  v(ldwl[296])
.save  v(ldwl[295])
.save  v(ldwl[294])
.save  v(ldwl[293])
.save  v(ldwl[292])
.save  v(ldwl[291])
.save  v(ldwl[290])
.save  v(ldwl[289])
.save  v(ldwl[288])
.save  v(ldwl[287])
.save  v(ldwl[286])
.save  v(ldwl[285])
.save  v(ldwl[284])
.save  v(ldwl[283])
.save  v(ldwl[282])
.save  v(ldwl[281])
.save  v(ldwl[280])
.save  v(ldwl[279])
.save  v(ldwl[278])
.save  v(ldwl[277])
.save  v(ldwl[276])
.save  v(ldwl[275])
.save  v(ldwl[274])
.save  v(ldwl[273])
.save  v(ldwl[272])
.save  v(ldwl[271])
.save  v(ldwl[270])
.save  v(ldwl[269])
.save  v(ldwl[268])
.save  v(ldwl[267])
.save  v(ldwl[266])
.save  v(ldwl[265])
.save  v(ldwl[264])
.save  v(ldwl[263])
.save  v(ldwl[262])
.save  v(ldwl[261])
.save  v(ldwl[260])
.save  v(ldwl[259])
.save  v(ldwl[258])
.save  v(ldwl[257])
.save  v(ldwl[256])
.save  v(ldwl[255])
.save  v(ldwl[254])
.save  v(ldwl[253])
.save  v(ldwl[252])
.save  v(ldwl[251])
.save  v(ldwl[250])
.save  v(ldwl[249])
.save  v(ldwl[248])
.save  v(ldwl[247])
.save  v(ldwl[246])
.save  v(ldwl[245])
.save  v(ldwl[244])
.save  v(ldwl[243])
.save  v(ldwl[242])
.save  v(ldwl[241])
.save  v(ldwl[240])
.save  v(ldwl[239])
.save  v(ldwl[238])
.save  v(ldwl[237])
.save  v(ldwl[236])
.save  v(ldwl[235])
.save  v(ldwl[234])
.save  v(ldwl[233])
.save  v(ldwl[232])
.save  v(ldwl[231])
.save  v(ldwl[230])
.save  v(ldwl[229])
.save  v(ldwl[228])
.save  v(ldwl[227])
.save  v(ldwl[226])
.save  v(ldwl[225])
.save  v(ldwl[224])
.save  v(ldwl[223])
.save  v(ldwl[222])
.save  v(ldwl[221])
.save  v(ldwl[220])
.save  v(ldwl[219])
.save  v(ldwl[218])
.save  v(ldwl[217])
.save  v(ldwl[216])
.save  v(ldwl[215])
.save  v(ldwl[214])
.save  v(ldwl[213])
.save  v(ldwl[212])
.save  v(ldwl[211])
.save  v(ldwl[210])
.save  v(ldwl[209])
.save  v(ldwl[208])
.save  v(ldwl[207])
.save  v(ldwl[206])
.save  v(ldwl[205])
.save  v(ldwl[204])
.save  v(ldwl[203])
.save  v(ldwl[202])
.save  v(ldwl[201])
.save  v(ldwl[200])
.save  v(ldwl[199])
.save  v(ldwl[198])
.save  v(ldwl[197])
.save  v(ldwl[196])
.save  v(ldwl[195])
.save  v(ldwl[194])
.save  v(ldwl[193])
.save  v(ldwl[192])
.save  v(ldwl[191])
.save  v(ldwl[190])
.save  v(ldwl[189])
.save  v(ldwl[188])
.save  v(ldwl[187])
.save  v(ldwl[186])
.save  v(ldwl[185])
.save  v(ldwl[184])
.save  v(ldwl[183])
.save  v(ldwl[182])
.save  v(ldwl[181])
.save  v(ldwl[180])
.save  v(ldwl[179])
.save  v(ldwl[178])
.save  v(ldwl[177])
.save  v(ldwl[176])
.save  v(ldwl[175])
.save  v(ldwl[174])
.save  v(ldwl[173])
.save  v(ldwl[172])
.save  v(ldwl[171])
.save  v(ldwl[170])
.save  v(ldwl[169])
.save  v(ldwl[168])
.save  v(ldwl[167])
.save  v(ldwl[166])
.save  v(ldwl[165])
.save  v(ldwl[164])
.save  v(ldwl[163])
.save  v(ldwl[162])
.save  v(ldwl[161])
.save  v(ldwl[160])
.save  v(ldwl[159])
.save  v(ldwl[158])
.save  v(ldwl[157])
.save  v(ldwl[156])
.save  v(ldwl[155])
.save  v(ldwl[154])
.save  v(ldwl[153])
.save  v(ldwl[152])
.save  v(ldwl[151])
.save  v(ldwl[150])
.save  v(ldwl[149])
.save  v(ldwl[148])
.save  v(ldwl[147])
.save  v(ldwl[146])
.save  v(ldwl[145])
.save  v(ldwl[144])
.save  v(ldwl[143])
.save  v(ldwl[142])
.save  v(ldwl[141])
.save  v(ldwl[140])
.save  v(ldwl[139])
.save  v(ldwl[138])
.save  v(ldwl[137])
.save  v(ldwl[136])
.save  v(ldwl[135])
.save  v(ldwl[134])
.save  v(ldwl[133])
.save  v(ldwl[132])
.save  v(ldwl[131])
.save  v(ldwl[130])
.save  v(ldwl[129])
.save  v(ldwl[128])
.save  v(ldwl[127])
.save  v(ldwl[126])
.save  v(ldwl[125])
.save  v(ldwl[124])
.save  v(ldwl[123])
.save  v(ldwl[122])
.save  v(ldwl[121])
.save  v(ldwl[120])
.save  v(ldwl[119])
.save  v(ldwl[118])
.save  v(ldwl[117])
.save  v(ldwl[116])
.save  v(ldwl[115])
.save  v(ldwl[114])
.save  v(ldwl[113])
.save  v(ldwl[112])
.save  v(ldwl[111])
.save  v(ldwl[110])
.save  v(ldwl[109])
.save  v(ldwl[108])
.save  v(ldwl[107])
.save  v(ldwl[106])
.save  v(ldwl[105])
.save  v(ldwl[104])
.save  v(ldwl[103])
.save  v(ldwl[102])
.save  v(ldwl[101])
.save  v(ldwl[100])
.save  v(ldwl[99])
.save  v(ldwl[98])
.save  v(ldwl[97])
.save  v(ldwl[96])
.save  v(ldwl[95])
.save  v(ldwl[94])
.save  v(ldwl[93])
.save  v(ldwl[92])
.save  v(ldwl[91])
.save  v(ldwl[90])
.save  v(ldwl[89])
.save  v(ldwl[88])
.save  v(ldwl[87])
.save  v(ldwl[86])
.save  v(ldwl[85])
.save  v(ldwl[84])
.save  v(ldwl[83])
.save  v(ldwl[82])
.save  v(ldwl[81])
.save  v(ldwl[80])
.save  v(ldwl[79])
.save  v(ldwl[78])
.save  v(ldwl[77])
.save  v(ldwl[76])
.save  v(ldwl[75])
.save  v(ldwl[74])
.save  v(ldwl[73])
.save  v(ldwl[72])
.save  v(ldwl[71])
.save  v(ldwl[70])
.save  v(ldwl[69])
.save  v(ldwl[68])
.save  v(ldwl[67])
.save  v(ldwl[66])
.save  v(ldwl[65])
.save  v(ldwl[64])
.save  v(ldwl[63])
.save  v(ldwl[62])
.save  v(ldwl[61])
.save  v(ldwl[60])
.save  v(ldwl[59])
.save  v(ldwl[58])
.save  v(ldwl[57])
.save  v(ldwl[56])
.save  v(ldwl[55])
.save  v(ldwl[54])
.save  v(ldwl[53])
.save  v(ldwl[52])
.save  v(ldwl[51])
.save  v(ldwl[50])
.save  v(ldwl[49])
.save  v(ldwl[48])
.save  v(ldwl[47])
.save  v(ldwl[46])
.save  v(ldwl[45])
.save  v(ldwl[44])
.save  v(ldwl[43])
.save  v(ldwl[42])
.save  v(ldwl[41])
.save  v(ldwl[40])
.save  v(ldwl[39])
.save  v(ldwl[38])
.save  v(ldwl[37])
.save  v(ldwl[36])
.save  v(ldwl[35])
.save  v(ldwl[34])
.save  v(ldwl[33])
.save  v(ldwl[32])
.save  v(ldwl[31])
.save  v(ldwl[30])
.save  v(ldwl[29])
.save  v(ldwl[28])
.save  v(ldwl[27])
.save  v(ldwl[26])
.save  v(ldwl[25])
.save  v(ldwl[24])
.save  v(ldwl[23])
.save  v(ldwl[22])
.save  v(ldwl[21])
.save  v(ldwl[20])
.save  v(ldwl[19])
.save  v(ldwl[18])
.save  v(ldwl[17])
.save  v(ldwl[16])
.save  v(ldwl[15])
.save  v(ldwl[14])
.save  v(ldwl[13])
.save  v(ldwl[12])
.save  v(ldwl[11])
.save  v(ldwl[10])
.save  v(ldwl[9])
.save  v(ldwl[8])
.save  v(ldwl[7])
.save  v(ldwl[6])
.save  v(ldwl[5])
.save  v(ldwl[4])
.save  v(ldwl[3])
.save  v(ldwl[2])
.save  v(ldwl[1])
.save  v(ldwl[0])
.save  v(ldbl[0])
.save  v(ldbl[16])
.save  v(ldbl[32])
.save  v(ldbl[1])
.save  v(ldbl[17])
.save  v(ldbl[33])
.save  v(ldbl[2])
.save  v(ldbl[18])
.save  v(ldbl[34])
**** begin user architecture code


.options SCALE=0.10
.param VCC=1.5
.temp 25
.param WPRECH=30u

vvss vss 0 0

** to generate following file:
** copy .../share/doc/xschem/rom8k/stimuli.rom8k to simulation directory
** then do 'Simulation->Utile Stimuli Editor (GUI)' and press 'Translate'
.include stimuli_rom8k.cir

* .op ALL  4n
*.dc vvcc 0 2 0.1
.save tran i(vvcc) i(vsa) i(vl) i(vdec)
.tran 0.2n 480n uic

** download models from here:
** http://www.amarketplaceofideas.com/wp-content/uploads/2014/11/180nm-V1.7z
** and save to 'models_rom8k.txt' in simulation directory
.include models_rom8k.txt



**** end user architecture code
**.ends

* expanding   symbol:  rom2_coldec.sym # of pins=4
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_coldec.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_coldec.sch
.subckt rom2_coldec  LDYMS LDY1[15] LDY1[14] LDY1[13] LDY1[12] LDY1[11] LDY1[10] LDY1[9] LDY1[8]
+ LDY1[7] LDY1[6] LDY1[5] LDY1[4] LDY1[3] LDY1[2] LDY1[1] LDY1[0] LDBL[15] LDBL[14] LDBL[13] LDBL[12]
+ LDBL[11] LDBL[10] LDBL[9] LDBL[8] LDBL[7] LDBL[6] LDBL[5] LDBL[4] LDBL[3] LDBL[2] LDBL[1] LDBL[0] VSS
*.opin LDYMS
*.ipin
*+ LDY1[15],LDY1[14],LDY1[13],LDY1[12],LDY1[11],LDY1[10],LDY1[9],LDY1[8],LDY1[7],LDY1[6],LDY1[5],LDY1[4],LDY1[3],LDY1[2],LDY1[1],LDY1[0]
*.ipin
*+ LDBL[15],LDBL[14],LDBL[13],LDBL[12],LDBL[11],LDBL[10],LDBL[9],LDBL[8],LDBL[7],LDBL[6],LDBL[5],LDBL[4],LDBL[3],LDBL[2],LDBL[1],LDBL[0]
*.ipin VSS
m96[15] LDBL[15] LDY1[15] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[14] LDBL[14] LDY1[14] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[13] LDBL[13] LDY1[13] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[12] LDBL[12] LDY1[12] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[11] LDBL[11] LDY1[11] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[10] LDBL[10] LDY1[10] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[9] LDBL[9] LDY1[9] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[8] LDBL[8] LDY1[8] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[7] LDBL[7] LDY1[7] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[6] LDBL[6] LDY1[6] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[5] LDBL[5] LDY1[5] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[4] LDBL[4] LDY1[4] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[3] LDBL[3] LDY1[3] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[2] LDBL[2] LDY1[2] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[1] LDBL[1] LDY1[1] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m96[0] LDBL[0] LDY1[0] LDYMS 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
c61 LDYMS VSS 20f m=1
.ends


* expanding   symbol:  rom2_sa.sym # of pins=8
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_sa.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_sa.sch
.subckt rom2_sa  LDQ LDCP LDYMS LDOE LDPRECH LDSAL vcc vss
*.opin LDQ
*.ipin LDCP
*.ipin LDYMS
*.ipin LDOE
*.ipin LDPRECH
*.ipin LDSAL
*.ipin vcc
*.ipin vss
x242 LDSALI LDSALI_B vcc vss lvnot wn=8.4u lln=2.4u wp=12u lp=2.4u m=1
x249 LDCP_B LDCP vcc vss lvnot wn=8.4u lln=2.4u wp=20u lp=2.4u m=1
x6 LDQ LDQIII LDOE vcc vss bts
x7 net1 LDQII LDSALI LDSALI_B vcc vss passhs WN=12u LN=1.2u WP=12u LP=1.2u
m6 LDQII LDQIB net2 0 cmosn w=24u l=2.4u ad='24u *4.4u' as='24u *4.4u' pd='24u *2 + 8.8u' ps='24u *2 + 8.8u'
+ m=1
m7 LDQII LDQIB net3 VCC cmosp w=24u l=2.4u ad='24u *4.4u' as='24u *4.4u' pd='24u *2 + 8.8u' ps='24u *2 + 8.8u'
+ m=1
m4 net2 LDSALI vss 0 cmosn w=24u l=2.4u ad='24u *4.4u' as='24u *4.4u' pd='24u *2 + 8.8u' ps='24u *2 + 8.8u'
+ m=1
m1 net3 LDSALI_B vcc VCC cmosp w=24u l=2.4u ad='24u *4.4u' as='24u *4.4u' pd='24u *2 + 8.8u' ps='24u *2 + 8.8u'
+ m=1
x8 net4 LDQII vcc vss lvnot wn=8.4u lln=2.4u wp=12u lp=2.4u m=1
x9 net1 net4 vcc vss lvnot wn=8.4u lln=2.4u wp=12u lp=2.4u m=1
c0 LDQII vss 3f m=1
c1 LDQIB vss 3f m=1
x228 LDQIII LDQII vcc vss lvnot wn=24u lln=2.4u wp=60u lp=2.4u m=1
x1 LDSALI_B LDSAL vcc vss lvnot wn=8.4u lln=2.4u wp=12u lp=2.4u m=1
xsacell LDCP_B LDPRECH vcc vss LDQI LDQIB LDYMS rom2_sacell
.save  v(ldqib)
.save  v(ldqii)
.save  v(ldcp_b)
.save  v(ldsali)
.save  v(ldqi)
.save  v(ldqiii)
.ends


* expanding   symbol:  rom2_addlatch.sym # of pins=7
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_addlatch.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_addlatch.sch
.subckt rom2_addlatch  LDEN_LAT LDAI[12] LDAI[11] LDAI[10] LDAI[9] LDAI[8] LDAI[7] LDAI[6] LDAI[5]
+ LDAI[4] LDAI[3] LDAI[2] LDAI[1] LDAI[0] LDEN LDCP_B LDA[12] LDA[11] LDA[10] LDA[9] LDA[8] LDA[7] LDA[6]
+ LDA[5] LDA[4] LDA[3] LDA[2] LDA[1] LDA[0] VCC VSS
*.opin LDEN_LAT
*.opin
*+ LDAI[12],LDAI[11],LDAI[10],LDAI[9],LDAI[8],LDAI[7],LDAI[6],LDAI[5],LDAI[4],LDAI[3],LDAI[2],LDAI[1],LDAI[0]
*.ipin LDEN
*.ipin LDCP_B
*.ipin LDA[12],LDA[11],LDA[10],LDA[9],LDA[8],LDA[7],LDA[6],LDA[5],LDA[4],LDA[3],LDA[2],LDA[1],LDA[0]
*.ipin VCC
*.ipin VSS
x0[12] LDA[12] LDCP_B VCC net1[12] VCC VSS VCC VSS LD2QHDX4stef
x0[11] LDA[11] LDCP_B VCC net1[11] VCC VSS VCC VSS LD2QHDX4stef
x0[10] LDA[10] LDCP_B VCC net1[10] VCC VSS VCC VSS LD2QHDX4stef
x0[9] LDA[9] LDCP_B VCC net1[9] VCC VSS VCC VSS LD2QHDX4stef
x0[8] LDA[8] LDCP_B VCC net1[8] VCC VSS VCC VSS LD2QHDX4stef
x0[7] LDA[7] LDCP_B VCC net1[7] VCC VSS VCC VSS LD2QHDX4stef
x0[6] LDA[6] LDCP_B VCC net1[6] VCC VSS VCC VSS LD2QHDX4stef
x0[5] LDA[5] LDCP_B VCC net1[5] VCC VSS VCC VSS LD2QHDX4stef
x0[4] LDA[4] LDCP_B VCC net1[4] VCC VSS VCC VSS LD2QHDX4stef
x0[3] LDA[3] LDCP_B VCC net1[3] VCC VSS VCC VSS LD2QHDX4stef
x0[2] LDA[2] LDCP_B VCC net1[2] VCC VSS VCC VSS LD2QHDX4stef
x0[1] LDA[1] LDCP_B VCC net1[1] VCC VSS VCC VSS LD2QHDX4stef
x0[0] LDA[0] LDCP_B VCC net1[0] VCC VSS VCC VSS LD2QHDX4stef
x9[12] LDAI[12] net2[12] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[11] LDAI[11] net2[11] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[10] LDAI[10] net2[10] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[9] LDAI[9] net2[9] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[8] LDAI[8] net2[8] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[7] LDAI[7] net2[7] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[6] LDAI[6] net2[6] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[5] LDAI[5] net2[5] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[4] LDAI[4] net2[4] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[3] LDAI[3] net2[3] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[2] LDAI[2] net2[2] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[1] LDAI[1] net2[1] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[0] LDAI[0] net2[0] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x10[12] net2[12] net1[12] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[11] net2[11] net1[11] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[10] net2[10] net1[10] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[9] net2[9] net1[9] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[8] net2[8] net1[8] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[7] net2[7] net1[7] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[6] net2[6] net1[6] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[5] net2[5] net1[5] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[4] net2[4] net1[4] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[3] net2[3] net1[3] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[2] net2[2] net1[2] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[1] net2[1] net1[1] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x10[0] net2[0] net1[0] vcc vss lvnot wn=16u lln=2.4u wp=40u lp=2.4u m=1
x3 LDEN LDCP_B VCC LDEN_LAT VCC VSS VCC VSS LD2QHDX4stef
x1[12] LDAI[12] net2[12] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[11] LDAI[11] net2[11] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[10] LDAI[10] net2[10] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[9] LDAI[9] net2[9] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[8] LDAI[8] net2[8] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[7] LDAI[7] net2[7] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[6] LDAI[6] net2[6] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[5] LDAI[5] net2[5] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[4] LDAI[4] net2[4] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[3] LDAI[3] net2[3] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[2] LDAI[2] net2[2] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[1] LDAI[1] net2[1] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x1[0] LDAI[0] net2[0] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
.ends


* expanding   symbol:  rom2_ctrl.sym # of pins=11
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_ctrl.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_ctrl.sch
.subckt rom2_ctrl  LDPRECH LDSAL LDCP_ROWDEC LDCP_SA LDCP_ADDLAT_B LDCP_COL_B LDEN_LAT LDCP VCC VSS
+ LDYMSREF
*.opin LDPRECH
*.opin LDSAL
*.opin LDCP_ROWDEC
*.opin LDCP_SA
*.opin LDCP_ADDLAT_B
*.opin LDCP_COL_B
*.ipin LDEN_LAT
*.ipin LDCP
*.ipin VCC
*.ipin VSS
*.iopin LDYMSREF
c84 LDCPB VSS 5f m=1
x392 LDCPB LDCP LDEN_LAT vcc vss lvnand2 wna=90u lna=2.4u wpa=60u lpa=2.4u wnb=90u lnb=2.4u wpb=60u
+ lpb=2.4u m=1
x394 LDCP_SA LDCPB vcc vss lvnot wn=8.4u lln=2.8u wp=40u lp=2.4u m=1
x395 LDCP_ROWDEC net3 vcc vss lvnot wn=15u lln=2.4u wp=40u lp=2.4u m=10
x396 net8 LDCPB vcc vss lvnot wn=15u lln=2.4u wp=40u lp=2.4u m=1
x397 net3 net8 vcc vss lvnot wn=15u lln=2.4u wp=40u lp=2.4u m=4
x405 LDCP_ADDLAT_B LDCP vcc vss lvnot wn=30u lln=2.4u wp=80u lp=2.4u m=1
x7 LDCP_REF_B VSS vcc vss lvnot wn=24u lln=2.4u wp=40u lp=2.4u m=1
x8 LDPRECHREF LDCPB LDOUTI VCC VSS lvnor2 wna=8.4u lna=2.4u wpa=70u lpa=2.4u wnb=8.4u lnb=2.4u
+ wpb=70u lpb=2.4u m=1
x18 net1 LDQ_B net2 VCC VSS lvnand2 wna=20u lna=2.4u wpa=36u lpa=2.4u wnb=20u lnb=2.4u wpb=36u
+ lpb=2.4u m=1
x3 net2 LDCP_REF net1 VCC VSS lvnand2 wna=30u lna=2.4u wpa=30u lpa=2.4u wnb=30u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
m15 net4 LDOUTI VSS 0 cmosn w=4u l=2.4u ad='4u *4.4u' as='4u *4.4u' pd='4u *2 + 8.8u' ps='4u *2 + 8.8u'
+ m=1
x25 net9 LDCP_REF LDQ_B LDOUTI VCC VSS lvnand3 wn=80u lln=2.4u wp=40u lp=2.4u m=1
x26 LDSAL net9 vcc vss lvnot wn=13u lln=2.4u wp=40u lp=2.4u m=4
x28 LDPRECH net10 vcc vss lvnot wn=13u lln=2.4u wp=40u lp=2.4u m=8
x4 LDCP_REF LDCPB vcc vss lvnot wn=13u lln=2.4u wp=40u lp=2.4u m=2
x1 LDCP_COL_B net11 vcc vss lvnot wn=20u lln=2.4u wp=44u lp=2.4u m=2
x6 net11 LDCPB vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x5 LDOUTIB net1 vcc vss lvnot wn=30u lln=2.4u wp=40u lp=2.4u m=1
x9 LDOUTI net2 vcc vss lvnot wn=12u lln=2.4u wp=30u lp=2.4u m=2
xsacell LDCPB LDPRECHREF VCC VSS LDQI LDQ_B LDYMSREF rom2_sacell
.save  v(ldcp_ref)
.save  v(ldprechref)
.save  v(ldouti)
.save  v(ldoutib)
.save  v(ldqi)
.save  v(ldq_b)
m1 net5 LDOUTI net4 0 cmosn w=4u l=2.4u ad='4u *4.4u' as='4u *4.4u' pd='4u *2 + 8.8u' ps='4u *2 + 8.8u'
+ m=1
x2 net10 LDOUTIB LDEN_LAT LDCP VCC VSS lvnand3 wn=80u lln=2.4u wp=60u lp=2.4u m=1
m2 net6 LDOUTI VSS 0 cmosn w=4u l=2.4u ad='4u *4.4u' as='4u *4.4u' pd='4u *2 + 8.8u' ps='4u *2 + 8.8u'
+ m=1
m0 net7 LDOUTI net6 0 cmosn w=4u l=2.4u ad='4u *4.4u' as='4u *4.4u' pd='4u *2 + 8.8u' ps='4u *2 + 8.8u'
+ m=1
.save  v(ldcpb)
.ends


* expanding   symbol:  rom2_predec3.sym # of pins=4
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_predec3.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_predec3.sch
.subckt rom2_predec3  LDZ[15] LDZ[14] LDZ[13] LDZ[12] LDZ[11] LDZ[10] LDZ[9] LDZ[8] LDZ[7] LDZ[6]
+ LDZ[5] LDZ[4] LDZ[3] LDZ[2] LDZ[1] LDZ[0] LDA[3] LDA[2] LDA[1] LDA[0] vcc vss
*.opin
*+ LDZ[15],LDZ[14],LDZ[13],LDZ[12],LDZ[11],LDZ[10],LDZ[9],LDZ[8],LDZ[7],LDZ[6],LDZ[5],LDZ[4],LDZ[3],LDZ[2],LDZ[1],LDZ[0]
*.ipin LDA[3],LDA[2],LDA[1],LDA[0]
*.ipin vcc
*.ipin vss
x325[15] net9[15] net10[15] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[14] net9[14] net10[14] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[13] net9[13] net10[13] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[12] net9[12] net10[12] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[11] net9[11] net10[11] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[10] net9[10] net10[10] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[9] net9[9] net10[9] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[8] net9[8] net10[8] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[7] net9[7] net10[7] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[6] net9[6] net10[6] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[5] net9[5] net10[5] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[4] net9[4] net10[4] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[3] net9[3] net10[3] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[2] net9[2] net10[2] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[1] net9[1] net10[1] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x325[0] net9[0] net10[0] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x8[15] LDZ[15] net9[15] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[14] LDZ[14] net9[14] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[13] LDZ[13] net9[13] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[12] LDZ[12] net9[12] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[11] LDZ[11] net9[11] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[10] LDZ[10] net9[10] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[9] LDZ[9] net9[9] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[8] LDZ[8] net9[8] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[7] LDZ[7] net9[7] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[6] LDZ[6] net9[6] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[5] LDZ[5] net9[5] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[4] LDZ[4] net9[4] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[3] LDZ[3] net9[3] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[2] LDZ[2] net9[2] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[1] LDZ[1] net9[1] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8[0] LDZ[0] net9[0] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9[15] net10[15] LDY[3] LDX[3] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[14] net10[14] LDY[3] LDX[2] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[13] net10[13] LDY[3] LDX[1] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[12] net10[12] LDY[3] LDX[0] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[11] net10[11] LDY[2] LDX[3] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[10] net10[10] LDY[2] LDX[2] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[9] net10[9] LDY[2] LDX[1] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[8] net10[8] LDY[2] LDX[0] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[7] net10[7] LDY[1] LDX[3] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[6] net10[6] LDY[1] LDX[2] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[5] net10[5] LDY[1] LDX[1] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[4] net10[4] LDY[1] LDX[0] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[3] net10[3] LDY[0] LDX[3] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[2] net10[2] LDY[0] LDX[2] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[1] net10[1] LDY[0] LDX[1] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[0] net10[0] LDY[0] LDX[0] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
c1[3] LDX[3] vss 14f m=1
c1[2] LDX[2] vss 14f m=1
c1[1] LDX[1] vss 14f m=1
c1[0] LDX[0] vss 14f m=1
c2[3] LDY[3] vss 14f m=1
c2[2] LDY[2] vss 14f m=1
c2[1] LDY[1] vss 14f m=1
c2[0] LDY[0] vss 14f m=1
x2 LDY[3] LDA[3] LDA[2] vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x3 LDY[2] LDA[3] net1 vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x4 LDY[1] net2 LDA[2] vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x6 LDY[0] net3 net4 vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x12 net1 LDA[2] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x1 net2 LDA[3] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x5 net4 LDA[2] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x7 net3 LDA[3] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x10 LDX[3] LDA[1] LDA[0] vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x20 LDX[2] LDA[1] net5 vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x11 LDX[1] net6 LDA[0] vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x13 LDX[0] net7 net8 vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x14 net5 LDA[0] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x15 net6 LDA[1] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x16 net8 LDA[0] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x17 net7 LDA[1] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x18[15] net9[15] net10[15] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[14] net9[14] net10[14] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[13] net9[13] net10[13] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[12] net9[12] net10[12] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[11] net9[11] net10[11] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[10] net9[10] net10[10] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[9] net9[9] net10[9] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[8] net9[8] net10[8] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[7] net9[7] net10[7] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[6] net9[6] net10[6] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[5] net9[5] net10[5] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[4] net9[4] net10[4] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[3] net9[3] net10[3] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[2] net9[2] net10[2] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[1] net9[1] net10[1] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x18[0] net9[0] net10[0] vcc vss lvnot wn=10u lln=2.4u wp=20u lp=2.4u m=1
x19[15] LDZ[15] net9[15] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[14] LDZ[14] net9[14] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[13] LDZ[13] net9[13] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[12] LDZ[12] net9[12] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[11] LDZ[11] net9[11] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[10] LDZ[10] net9[10] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[9] LDZ[9] net9[9] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[8] LDZ[8] net9[8] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[7] LDZ[7] net9[7] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[6] LDZ[6] net9[6] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[5] LDZ[5] net9[5] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[4] LDZ[4] net9[4] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[3] LDZ[3] net9[3] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[2] LDZ[2] net9[2] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[1] LDZ[1] net9[1] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x19[0] LDZ[0] net9[0] vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
.ends


* expanding   symbol:  rom3_rowdec.sym # of pins=7
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom3_rowdec.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom3_rowdec.sch
.subckt rom3_rowdec  LDWL[15] LDWL[14] LDWL[13] LDWL[12] LDWL[11] LDWL[10] LDWL[9] LDWL[8] LDWL[7]
+ LDWL[6] LDWL[5] LDWL[4] LDWL[3] LDWL[2] LDWL[1] LDWL[0] LDL1X[15] LDL1X[14] LDL1X[13] LDL1X[12] LDL1X[11]
+ LDL1X[10] LDL1X[9] LDL1X[8] LDL1X[7] LDL1X[6] LDL1X[5] LDL1X[4] LDL1X[3] LDL1X[2] LDL1X[1] LDL1X[0] LDL2X
+ LDL3X LDCP VSS VCC
*.opin
*+ LDWL[15],LDWL[14],LDWL[13],LDWL[12],LDWL[11],LDWL[10],LDWL[9],LDWL[8],LDWL[7],LDWL[6],LDWL[5],LDWL[4],LDWL[3],LDWL[2],LDWL[1],LDWL[0]
*.ipin
*+ LDL1X[15],LDL1X[14],LDL1X[13],LDL1X[12],LDL1X[11],LDL1X[10],LDL1X[9],LDL1X[8],LDL1X[7],LDL1X[6],LDL1X[5],LDL1X[4],LDL1X[3],LDL1X[2],LDL1X[1],LDL1X[0]
*.ipin LDL2X
*.ipin LDL3X
*.ipin LDCP
*.ipin VSS
*.ipin VCC
m0[15] net1[15] LDL1X[15] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u'
+ ps='14u *2 + 8.8u' m=1
m0[14] net1[14] LDL1X[14] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u'
+ ps='14u *2 + 8.8u' m=1
m0[13] net1[13] LDL1X[13] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u'
+ ps='14u *2 + 8.8u' m=1
m0[12] net1[12] LDL1X[12] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u'
+ ps='14u *2 + 8.8u' m=1
m0[11] net1[11] LDL1X[11] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u'
+ ps='14u *2 + 8.8u' m=1
m0[10] net1[10] LDL1X[10] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u'
+ ps='14u *2 + 8.8u' m=1
m0[9] net1[9] LDL1X[9] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[8] net1[8] LDL1X[8] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[7] net1[7] LDL1X[7] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[6] net1[6] LDL1X[6] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[5] net1[5] LDL1X[5] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[4] net1[4] LDL1X[4] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[3] net1[3] LDL1X[3] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[2] net1[2] LDL1X[2] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[1] net1[1] LDL1X[1] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
m0[0] net1[0] LDL1X[0] LDL1X_S 0 cmosn w=14u l=2u ad='14u *4.4u' as='14u *4.4u' pd='14u *2 + 8.8u' ps='14u *2 + 8.8u'
+ m=1
c1[15] LDWL_B[15] VSS 3f m=1
c1[14] LDWL_B[14] VSS 3f m=1
c1[13] LDWL_B[13] VSS 3f m=1
c1[12] LDWL_B[12] VSS 3f m=1
c1[11] LDWL_B[11] VSS 3f m=1
c1[10] LDWL_B[10] VSS 3f m=1
c1[9] LDWL_B[9] VSS 3f m=1
c1[8] LDWL_B[8] VSS 3f m=1
c1[7] LDWL_B[7] VSS 3f m=1
c1[6] LDWL_B[6] VSS 3f m=1
c1[5] LDWL_B[5] VSS 3f m=1
c1[4] LDWL_B[4] VSS 3f m=1
c1[3] LDWL_B[3] VSS 3f m=1
c1[2] LDWL_B[2] VSS 3f m=1
c1[1] LDWL_B[1] VSS 3f m=1
c1[0] LDWL_B[0] VSS 3f m=1
x2[15] LDWL[15] LDWL_B[15] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[14] LDWL[14] LDWL_B[14] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[13] LDWL[13] LDWL_B[13] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[12] LDWL[12] LDWL_B[12] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[11] LDWL[11] LDWL_B[11] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[10] LDWL[10] LDWL_B[10] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[9] LDWL[9] LDWL_B[9] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[8] LDWL[8] LDWL_B[8] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[7] LDWL[7] LDWL_B[7] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[6] LDWL[6] LDWL_B[6] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[5] LDWL[5] LDWL_B[5] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[4] LDWL[4] LDWL_B[4] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[3] LDWL[3] LDWL_B[3] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[2] LDWL[2] LDWL_B[2] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[1] LDWL[1] LDWL_B[1] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
x2[0] LDWL[0] LDWL_B[0] vcc vss lvnot wn=24u lln=2.4u wp=120u lp=2.4u m=1
m3[15] LDWL_B[15] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u'
+ ps='8.4u *2 + 8.8u' m=1
m3[14] LDWL_B[14] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u'
+ ps='8.4u *2 + 8.8u' m=1
m3[13] LDWL_B[13] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u'
+ ps='8.4u *2 + 8.8u' m=1
m3[12] LDWL_B[12] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u'
+ ps='8.4u *2 + 8.8u' m=1
m3[11] LDWL_B[11] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u'
+ ps='8.4u *2 + 8.8u' m=1
m3[10] LDWL_B[10] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u'
+ ps='8.4u *2 + 8.8u' m=1
m3[9] LDWL_B[9] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[8] LDWL_B[8] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[7] LDWL_B[7] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[6] LDWL_B[6] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[5] LDWL_B[5] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[4] LDWL_B[4] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[3] LDWL_B[3] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[2] LDWL_B[2] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[1] LDWL_B[1] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m3[0] LDWL_B[0] VSS VCC VCC cmosp w=8.4u l=8.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m4[15] LDWL_B[15] LDCP net1[15] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u'
+ ps='19u *2 + 8.8u' m=1
m4[14] LDWL_B[14] LDCP net1[14] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u'
+ ps='19u *2 + 8.8u' m=1
m4[13] LDWL_B[13] LDCP net1[13] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u'
+ ps='19u *2 + 8.8u' m=1
m4[12] LDWL_B[12] LDCP net1[12] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u'
+ ps='19u *2 + 8.8u' m=1
m4[11] LDWL_B[11] LDCP net1[11] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u'
+ ps='19u *2 + 8.8u' m=1
m4[10] LDWL_B[10] LDCP net1[10] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u'
+ ps='19u *2 + 8.8u' m=1
m4[9] LDWL_B[9] LDCP net1[9] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[8] LDWL_B[8] LDCP net1[8] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[7] LDWL_B[7] LDCP net1[7] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[6] LDWL_B[6] LDCP net1[6] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[5] LDWL_B[5] LDCP net1[5] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[4] LDWL_B[4] LDCP net1[4] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[3] LDWL_B[3] LDCP net1[3] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[2] LDWL_B[2] LDCP net1[2] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[1] LDWL_B[1] LDCP net1[1] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m4[0] LDWL_B[0] LDCP net1[0] 0 cmosn w=19u l=2.4u ad='19u *4.4u' as='19u *4.4u' pd='19u *2 + 8.8u' ps='19u *2 + 8.8u'
+ m=1
m1 net2 LDL3X VSS 0 cmosn w=40u l=2.4u ad='40u *4.4u' as='40u *4.4u' pd='40u *2 + 8.8u' ps='40u *2 + 8.8u'
+ m=1
m2 LDL1X_S LDL2X net2 0 cmosn w=40u l=2.4u ad='40u *4.4u' as='40u *4.4u' pd='40u *2 + 8.8u' ps='40u *2 + 8.8u'
+ m=1
m5 LDL1X_S LDL2X VCC VCC cmosp w=8.4u l=2.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
m6 LDL1X_S LDL3X VCC VCC cmosp w=8.4u l=2.4u ad='8.4u *4.4u' as='8.4u *4.4u' pd='8.4u *2 + 8.8u' ps='8.4u *2 + 8.8u'
+ m=1
.ends


* expanding   symbol:  rom2_predec1.sym # of pins=4
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_predec1.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_predec1.sch
.subckt rom2_predec1  LDZ[15] LDZ[14] LDZ[13] LDZ[12] LDZ[11] LDZ[10] LDZ[9] LDZ[8] LDZ[7] LDZ[6]
+ LDZ[5] LDZ[4] LDZ[3] LDZ[2] LDZ[1] LDZ[0] LDA[3] LDA[2] LDA[1] LDA[0] vcc vss
*.opin
*+ LDZ[15],LDZ[14],LDZ[13],LDZ[12],LDZ[11],LDZ[10],LDZ[9],LDZ[8],LDZ[7],LDZ[6],LDZ[5],LDZ[4],LDZ[3],LDZ[2],LDZ[1],LDZ[0]
*.ipin LDA[3],LDA[2],LDA[1],LDA[0]
*.ipin vcc
*.ipin vss
x325[15] net9[15] LDZI[15] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[14] net9[14] LDZI[14] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[13] net9[13] LDZI[13] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[12] net9[12] LDZI[12] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[11] net9[11] LDZI[11] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[10] net9[10] LDZI[10] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[9] net9[9] LDZI[9] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[8] net9[8] LDZI[8] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[7] net9[7] LDZI[7] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[6] net9[6] LDZI[6] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[5] net9[5] LDZI[5] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[4] net9[4] LDZI[4] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[3] net9[3] LDZI[3] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[2] net9[2] LDZI[2] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[1] net9[1] LDZI[1] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x325[0] net9[0] LDZI[0] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x8[15] LDZ[15] net9[15] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[14] LDZ[14] net9[14] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[13] LDZ[13] net9[13] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[12] LDZ[12] net9[12] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[11] LDZ[11] net9[11] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[10] LDZ[10] net9[10] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[9] LDZ[9] net9[9] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[8] LDZ[8] net9[8] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[7] LDZ[7] net9[7] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[6] LDZ[6] net9[6] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[5] LDZ[5] net9[5] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[4] LDZ[4] net9[4] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[3] LDZ[3] net9[3] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[2] LDZ[2] net9[2] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[1] LDZ[1] net9[1] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x8[0] LDZ[0] net9[0] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x9[15] LDZI[15] LDY[3] LDX[3] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[14] LDZI[14] LDY[3] LDX[2] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[13] LDZI[13] LDY[3] LDX[1] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[12] LDZI[12] LDY[3] LDX[0] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[11] LDZI[11] LDY[2] LDX[3] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[10] LDZI[10] LDY[2] LDX[2] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[9] LDZI[9] LDY[2] LDX[1] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[8] LDZI[8] LDY[2] LDX[0] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[7] LDZI[7] LDY[1] LDX[3] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[6] LDZI[6] LDY[1] LDX[2] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[5] LDZI[5] LDY[1] LDX[1] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[4] LDZI[4] LDY[1] LDX[0] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[3] LDZI[3] LDY[0] LDX[3] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[2] LDZI[2] LDY[0] LDX[2] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[1] LDZI[1] LDY[0] LDX[1] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
x9[0] LDZI[0] LDY[0] LDX[0] vcc vss lvnor2 wna=10u lna=2.4u wpa=40u lpa=2.4u wnb=10u lnb=2.4u
+ wpb=40u lpb=2.4u m=1
c1[3] LDX[3] vss 35f m=1
c1[2] LDX[2] vss 35f m=1
c1[1] LDX[1] vss 35f m=1
c1[0] LDX[0] vss 35f m=1
c2[3] LDY[3] vss 16f m=1
c2[2] LDY[2] vss 16f m=1
c2[1] LDY[1] vss 16f m=1
c2[0] LDY[0] vss 16f m=1
x2 LDY[3] LDA[3] LDA[2] vcc vss lvnand2 wna=20u lna=2.4u wpa=30u lpa=2.4u wnb=20u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
x3 LDY[2] LDA[3] net1 vcc vss lvnand2 wna=20u lna=2.4u wpa=30u lpa=2.4u wnb=20u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
x4 LDY[1] net2 LDA[2] vcc vss lvnand2 wna=20u lna=2.4u wpa=30u lpa=2.4u wnb=20u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
x6 LDY[0] net3 net4 vcc vss lvnand2 wna=20u lna=2.4u wpa=30u lpa=2.4u wnb=20u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
x12 net1 LDA[2] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x1 net2 LDA[3] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x5 net4 LDA[2] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x7 net3 LDA[3] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x10 LDX[3] LDA[1] LDA[0] vcc vss lvnand2 wna=20u lna=2.4u wpa=30u lpa=2.4u wnb=20u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
x20 LDX[2] LDA[1] net5 vcc vss lvnand2 wna=20u lna=2.4u wpa=30u lpa=2.4u wnb=20u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
x11 LDX[1] net6 LDA[0] vcc vss lvnand2 wna=20u lna=2.4u wpa=30u lpa=2.4u wnb=20u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
x13 LDX[0] net7 net8 vcc vss lvnand2 wna=20u lna=2.4u wpa=30u lpa=2.4u wnb=20u lnb=2.4u wpb=30u
+ lpb=2.4u m=1
x14 net5 LDA[0] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x15 net6 LDA[1] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x16 net8 LDA[0] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x17 net7 LDA[1] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x18[15] net9[15] LDZI[15] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[14] net9[14] LDZI[14] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[13] net9[13] LDZI[13] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[12] net9[12] LDZI[12] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[11] net9[11] LDZI[11] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[10] net9[10] LDZI[10] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[9] net9[9] LDZI[9] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[8] net9[8] LDZI[8] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[7] net9[7] LDZI[7] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[6] net9[6] LDZI[6] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[5] net9[5] LDZI[5] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[4] net9[4] LDZI[4] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[3] net9[3] LDZI[3] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[2] net9[2] LDZI[2] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[1] net9[1] LDZI[1] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x18[0] net9[0] LDZI[0] vcc vss lvnot wn=20u lln=2.4u wp=40u lp=2.4u m=1
x19[15] LDZ[15] net9[15] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[14] LDZ[14] net9[14] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[13] LDZ[13] net9[13] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[12] LDZ[12] net9[12] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[11] LDZ[11] net9[11] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[10] LDZ[10] net9[10] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[9] LDZ[9] net9[9] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[8] LDZ[8] net9[8] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[7] LDZ[7] net9[7] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[6] LDZ[6] net9[6] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[5] LDZ[5] net9[5] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[4] LDZ[4] net9[4] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[3] LDZ[3] net9[3] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[2] LDZ[2] net9[2] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[1] LDZ[1] net9[1] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x19[0] LDZ[0] net9[0] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[15] LDZ[15] net9[15] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[14] LDZ[14] net9[14] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[13] LDZ[13] net9[13] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[12] LDZ[12] net9[12] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[11] LDZ[11] net9[11] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[10] LDZ[10] net9[10] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[9] LDZ[9] net9[9] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[8] LDZ[8] net9[8] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[7] LDZ[7] net9[7] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[6] LDZ[6] net9[6] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[5] LDZ[5] net9[5] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[4] LDZ[4] net9[4] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[3] LDZ[3] net9[3] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[2] LDZ[2] net9[2] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[1] LDZ[1] net9[1] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x21[0] LDZ[0] net9[0] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[15] LDZ[15] net9[15] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[14] LDZ[14] net9[14] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[13] LDZ[13] net9[13] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[12] LDZ[12] net9[12] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[11] LDZ[11] net9[11] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[10] LDZ[10] net9[10] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[9] LDZ[9] net9[9] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[8] LDZ[8] net9[8] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[7] LDZ[7] net9[7] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[6] LDZ[6] net9[6] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[5] LDZ[5] net9[5] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[4] LDZ[4] net9[4] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[3] LDZ[3] net9[3] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[2] LDZ[2] net9[2] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[1] LDZ[1] net9[1] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
x22[0] LDZ[0] net9[0] vcc vss lvnot wn=30u lln=2.4u wp=60u lp=2.4u m=1
.ends


* expanding   symbol:  rom2_predec4.sym # of pins=5
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_predec4.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_predec4.sch
.subckt rom2_predec4  LDA[4] LDA[3] LDA[2] LDA[1] LDA[0] vcc vss LDL2X[3] LDL2X[2] LDL2X[1] LDL2X[0]
+ LDL3X[7] LDL3X[6] LDL3X[5] LDL3X[4] LDL3X[3] LDL3X[2] LDL3X[1] LDL3X[0]
*.ipin LDA[4],LDA[3],LDA[2],LDA[1],LDA[0]
*.ipin vcc
*.ipin vss
*.opin LDL2X[3],LDL2X[2],LDL2X[1],LDL2X[0]
*.opin LDL3X[7],LDL3X[6],LDL3X[5],LDL3X[4],LDL3X[3],LDL3X[2],LDL3X[1],LDL3X[0]
x10 net17 LDA[1] LDA[0] vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x2 net18 LDA[1] net1 vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x11 net19 net2 LDA[0] vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x13 net20 net3 net4 vcc vss lvnand2 wna=20u lna=2.4u wpa=20u lpa=2.4u wnb=20u lnb=2.4u wpb=20u
+ lpb=2.4u m=1
x17 net1 LDA[0] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x18 net2 LDA[1] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x19 net4 LDA[0] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x20 net3 LDA[1] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x5 net21 LDA[4] LDA[3] LDA[2] vcc vss lvnand3 wn=30u lln=2.4u wp=20u lp=2.4u m=1
x6 LDL3X[7] net21 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x14 net22 LDA[4] LDA[3] net5 vcc vss lvnand3 wn=30u lln=2.4u wp=20u lp=2.4u m=1
x15 LDL3X[6] net22 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x22 net5 LDA[2] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x23 net23 LDA[4] net6 LDA[2] vcc vss lvnand3 wn=30u lln=2.4u wp=20u lp=2.4u m=1
x24 LDL2X[3] net17 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x26 net6 LDA[3] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x28 net24 LDA[4] net7 net8 vcc vss lvnand3 wn=30u lln=2.4u wp=20u lp=2.4u m=1
x29 LDL3X[4] net24 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x31 net7 LDA[3] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x32 net8 LDA[2] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x33 net25 net9 LDA[3] LDA[2] vcc vss lvnand3 wn=30u lln=2.4u wp=20u lp=2.4u m=1
x34 LDL3X[3] net25 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x35 net9 LDA[4] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x38 net26 net11 LDA[3] net10 vcc vss lvnand3 wn=30u lln=2.4u wp=20u lp=2.4u m=1
x39 LDL3X[2] net26 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x40 net11 LDA[4] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x42 net10 LDA[2] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x43 net27 net13 net12 LDA[2] vcc vss lvnand3 wn=30u lln=2.4u wp=20u lp=2.4u m=1
x44 LDL3X[1] net27 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x45 net13 LDA[4] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x46 net12 LDA[3] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x48 net28 net16 net14 net15 vcc vss lvnand3 wn=30u lln=2.4u wp=20u lp=2.4u m=1
x49 LDL3X[0] net28 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x50 net16 LDA[4] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x51 net14 LDA[3] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x52 net15 LDA[2] vcc vss lvnot wn=8.4u lln=2.4u wp=16u lp=2.4u m=1
x1 LDL2X[2] net18 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x3 LDL2X[1] net19 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x0 LDL2X[0] net20 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x4 LDL3X[5] net23 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x7 LDL3X[7] net21 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x8 LDL3X[6] net22 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x9 LDL2X[3] net17 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x12 LDL3X[4] net24 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x16 LDL3X[3] net25 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x21 LDL3X[2] net26 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x25 LDL3X[1] net27 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x27 LDL3X[0] net28 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x30 LDL2X[2] net18 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x36 LDL2X[1] net19 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x37 LDL2X[0] net20 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
x41 LDL3X[5] net23 vcc vss lvnot wn=24u lln=2.4u wp=80u lp=2.4u m=1
.ends


* expanding   symbol:  rom2_coldec_ref.sym # of pins=4
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_coldec_ref.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_coldec_ref.sch
.subckt rom2_coldec_ref  LDYMSREF LDBLREF VCC VSS
*.opin LDYMSREF
*.ipin LDBLREF
*.ipin VCC
*.ipin VSS
m1 LDBLREF VCC LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
c61 LDYMSREF VSS 20f m=1
m2[15] net1[14] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[14] net1[13] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[13] net1[12] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[12] net1[11] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[11] net1[10] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[10] net1[9] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[9] net1[8] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[8] net1[7] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[7] net1[6] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[6] net1[5] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[5] net1[4] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[4] net1[3] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[3] net1[2] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[2] net1[1] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
m2[1] net1[0] VSS LDYMSREF 0 cmosn w=50u l=2u ad='50u *4.4u' as='50u *4.4u' pd='50u *2 + 8.8u' ps='50u *2 + 8.8u'
+ m=1
.ends


* expanding   symbol:  rom3_array_ref.sym # of pins=3
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom3_array_ref.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom3_array_ref.sch
.subckt rom3_array_ref  LDWL[511] LDWL[510] LDWL[509] LDWL[508] LDWL[507] LDWL[506] LDWL[505]
+ LDWL[504] LDWL[503] LDWL[502] LDWL[501] LDWL[500] LDWL[499] LDWL[498] LDWL[497] LDWL[496] LDWL[495] LDWL[494]
+ LDWL[493] LDWL[492] LDWL[491] LDWL[490] LDWL[489] LDWL[488] LDWL[487] LDWL[486] LDWL[485] LDWL[484] LDWL[483]
+ LDWL[482] LDWL[481] LDWL[480] LDWL[479] LDWL[478] LDWL[477] LDWL[476] LDWL[475] LDWL[474] LDWL[473] LDWL[472]
+ LDWL[471] LDWL[470] LDWL[469] LDWL[468] LDWL[467] LDWL[466] LDWL[465] LDWL[464] LDWL[463] LDWL[462] LDWL[461]
+ LDWL[460] LDWL[459] LDWL[458] LDWL[457] LDWL[456] LDWL[455] LDWL[454] LDWL[453] LDWL[452] LDWL[451] LDWL[450]
+ LDWL[449] LDWL[448] LDWL[447] LDWL[446] LDWL[445] LDWL[444] LDWL[443] LDWL[442] LDWL[441] LDWL[440] LDWL[439]
+ LDWL[438] LDWL[437] LDWL[436] LDWL[435] LDWL[434] LDWL[433] LDWL[432] LDWL[431] LDWL[430] LDWL[429] LDWL[428]
+ LDWL[427] LDWL[426] LDWL[425] LDWL[424] LDWL[423] LDWL[422] LDWL[421] LDWL[420] LDWL[419] LDWL[418] LDWL[417]
+ LDWL[416] LDWL[415] LDWL[414] LDWL[413] LDWL[412] LDWL[411] LDWL[410] LDWL[409] LDWL[408] LDWL[407] LDWL[406]
+ LDWL[405] LDWL[404] LDWL[403] LDWL[402] LDWL[401] LDWL[400] LDWL[399] LDWL[398] LDWL[397] LDWL[396] LDWL[395]
+ LDWL[394] LDWL[393] LDWL[392] LDWL[391] LDWL[390] LDWL[389] LDWL[388] LDWL[387] LDWL[386] LDWL[385] LDWL[384]
+ LDWL[383] LDWL[382] LDWL[381] LDWL[380] LDWL[379] LDWL[378] LDWL[377] LDWL[376] LDWL[375] LDWL[374] LDWL[373]
+ LDWL[372] LDWL[371] LDWL[370] LDWL[369] LDWL[368] LDWL[367] LDWL[366] LDWL[365] LDWL[364] LDWL[363] LDWL[362]
+ LDWL[361] LDWL[360] LDWL[359] LDWL[358] LDWL[357] LDWL[356] LDWL[355] LDWL[354] LDWL[353] LDWL[352] LDWL[351]
+ LDWL[350] LDWL[349] LDWL[348] LDWL[347] LDWL[346] LDWL[345] LDWL[344] LDWL[343] LDWL[342] LDWL[341] LDWL[340]
+ LDWL[339] LDWL[338] LDWL[337] LDWL[336] LDWL[335] LDWL[334] LDWL[333] LDWL[332] LDWL[331] LDWL[330] LDWL[329]
+ LDWL[328] LDWL[327] LDWL[326] LDWL[325] LDWL[324] LDWL[323] LDWL[322] LDWL[321] LDWL[320] LDWL[319] LDWL[318]
+ LDWL[317] LDWL[316] LDWL[315] LDWL[314] LDWL[313] LDWL[312] LDWL[311] LDWL[310] LDWL[309] LDWL[308] LDWL[307]
+ LDWL[306] LDWL[305] LDWL[304] LDWL[303] LDWL[302] LDWL[301] LDWL[300] LDWL[299] LDWL[298] LDWL[297] LDWL[296]
+ LDWL[295] LDWL[294] LDWL[293] LDWL[292] LDWL[291] LDWL[290] LDWL[289] LDWL[288] LDWL[287] LDWL[286] LDWL[285]
+ LDWL[284] LDWL[283] LDWL[282] LDWL[281] LDWL[280] LDWL[279] LDWL[278] LDWL[277] LDWL[276] LDWL[275] LDWL[274]
+ LDWL[273] LDWL[272] LDWL[271] LDWL[270] LDWL[269] LDWL[268] LDWL[267] LDWL[266] LDWL[265] LDWL[264] LDWL[263]
+ LDWL[262] LDWL[261] LDWL[260] LDWL[259] LDWL[258] LDWL[257] LDWL[256] LDWL[255] LDWL[254] LDWL[253] LDWL[252]
+ LDWL[251] LDWL[250] LDWL[249] LDWL[248] LDWL[247] LDWL[246] LDWL[245] LDWL[244] LDWL[243] LDWL[242] LDWL[241]
+ LDWL[240] LDWL[239] LDWL[238] LDWL[237] LDWL[236] LDWL[235] LDWL[234] LDWL[233] LDWL[232] LDWL[231] LDWL[230]
+ LDWL[229] LDWL[228] LDWL[227] LDWL[226] LDWL[225] LDWL[224] LDWL[223] LDWL[222] LDWL[221] LDWL[220] LDWL[219]
+ LDWL[218] LDWL[217] LDWL[216] LDWL[215] LDWL[214] LDWL[213] LDWL[212] LDWL[211] LDWL[210] LDWL[209] LDWL[208]
+ LDWL[207] LDWL[206] LDWL[205] LDWL[204] LDWL[203] LDWL[202] LDWL[201] LDWL[200] LDWL[199] LDWL[198] LDWL[197]
+ LDWL[196] LDWL[195] LDWL[194] LDWL[193] LDWL[192] LDWL[191] LDWL[190] LDWL[189] LDWL[188] LDWL[187] LDWL[186]
+ LDWL[185] LDWL[184] LDWL[183] LDWL[182] LDWL[181] LDWL[180] LDWL[179] LDWL[178] LDWL[177] LDWL[176] LDWL[175]
+ LDWL[174] LDWL[173] LDWL[172] LDWL[171] LDWL[170] LDWL[169] LDWL[168] LDWL[167] LDWL[166] LDWL[165] LDWL[164]
+ LDWL[163] LDWL[162] LDWL[161] LDWL[160] LDWL[159] LDWL[158] LDWL[157] LDWL[156] LDWL[155] LDWL[154] LDWL[153]
+ LDWL[152] LDWL[151] LDWL[150] LDWL[149] LDWL[148] LDWL[147] LDWL[146] LDWL[145] LDWL[144] LDWL[143] LDWL[142]
+ LDWL[141] LDWL[140] LDWL[139] LDWL[138] LDWL[137] LDWL[136] LDWL[135] LDWL[134] LDWL[133] LDWL[132] LDWL[131]
+ LDWL[130] LDWL[129] LDWL[128] LDWL[127] LDWL[126] LDWL[125] LDWL[124] LDWL[123] LDWL[122] LDWL[121] LDWL[120]
+ LDWL[119] LDWL[118] LDWL[117] LDWL[116] LDWL[115] LDWL[114] LDWL[113] LDWL[112] LDWL[111] LDWL[110] LDWL[109]
+ LDWL[108] LDWL[107] LDWL[106] LDWL[105] LDWL[104] LDWL[103] LDWL[102] LDWL[101] LDWL[100] LDWL[99] LDWL[98]
+ LDWL[97] LDWL[96] LDWL[95] LDWL[94] LDWL[93] LDWL[92] LDWL[91] LDWL[90] LDWL[89] LDWL[88] LDWL[87] LDWL[86]
+ LDWL[85] LDWL[84] LDWL[83] LDWL[82] LDWL[81] LDWL[80] LDWL[79] LDWL[78] LDWL[77] LDWL[76] LDWL[75] LDWL[74]
+ LDWL[73] LDWL[72] LDWL[71] LDWL[70] LDWL[69] LDWL[68] LDWL[67] LDWL[66] LDWL[65] LDWL[64] LDWL[63] LDWL[62]
+ LDWL[61] LDWL[60] LDWL[59] LDWL[58] LDWL[57] LDWL[56] LDWL[55] LDWL[54] LDWL[53] LDWL[52] LDWL[51] LDWL[50]
+ LDWL[49] LDWL[48] LDWL[47] LDWL[46] LDWL[45] LDWL[44] LDWL[43] LDWL[42] LDWL[41] LDWL[40] LDWL[39] LDWL[38]
+ LDWL[37] LDWL[36] LDWL[35] LDWL[34] LDWL[33] LDWL[32] LDWL[31] LDWL[30] LDWL[29] LDWL[28] LDWL[27] LDWL[26]
+ LDWL[25] LDWL[24] LDWL[23] LDWL[22] LDWL[21] LDWL[20] LDWL[19] LDWL[18] LDWL[17] LDWL[16] LDWL[15] LDWL[14]
+ LDWL[13] LDWL[12] LDWL[11] LDWL[10] LDWL[9] LDWL[8] LDWL[7] LDWL[6] LDWL[5] LDWL[4] LDWL[3] LDWL[2] LDWL[1]
+ LDWL[0] vss LDBLREF
*.ipin
*+ LDWL[511],LDWL[510],LDWL[509],LDWL[508],LDWL[507],LDWL[506],LDWL[505],LDWL[504],LDWL[503],LDWL[502],LDWL[501],LDWL[500],LDWL[499],LDWL[498],LDWL[497],LDWL[496],LDWL[495],LDWL[494],LDWL[493],LDWL[492],LDWL[491],LDWL[490],LDWL[489],LDWL[488],LDWL[487],LDWL[486],LDWL[485],LDWL[484],LDWL[483],LDWL[482],LDWL[481],LDWL[480],LDWL[479],LDWL[478],LDWL[477],LDWL[476],LDWL[475],LDWL[474],LDWL[473],LDWL[472],LDWL[471],LDWL[470],LDWL[469],LDWL[468],LDWL[467],LDWL[466],LDWL[465],LDWL[464],LDWL[463],LDWL[462],LDWL[461],LDWL[460],LDWL[459],LDWL[458],LDWL[457],LDWL[456],LDWL[455],LDWL[454],LDWL[453],LDWL[452],LDWL[451],LDWL[450],LDWL[449],LDWL[448],LDWL[447],LDWL[446],LDWL[445],LDWL[444],LDWL[443],LDWL[442],LDWL[441],LDWL[440],LDWL[439],LDWL[438],LDWL[437],LDWL[436],LDWL[435],LDWL[434],LDWL[433],LDWL[432],LDWL[431],LDWL[430],LDWL[429],LDWL[428],LDWL[427],LDWL[426],LDWL[425],LDWL[424],LDWL[423],LDWL[422],LDWL[421],LDWL[420],LDWL[419],LDWL[418],LDWL[417],LDWL[416],LDWL[415],LDWL[414],LDWL[413],LDWL[412],LDWL[411],LDWL[410],LDWL[409],LDWL[408],LDWL[407],LDWL[406],LDWL[405],LDWL[404],LDWL[403],LDWL[402],LDWL[401],LDWL[400],LDWL[399],LDWL[398],LDWL[397],LDWL[396],LDWL[395],LDWL[394],LDWL[393],LDWL[392],LDWL[391],LDWL[390],LDWL[389],LDWL[388],LDWL[387],LDWL[386],LDWL[385],LDWL[384],LDWL[383],LDWL[382],LDWL[381],LDWL[380],LDWL[379],LDWL[378],LDWL[377],LDWL[376],LDWL[375],LDWL[374],LDWL[373],LDWL[372],LDWL[371],LDWL[370],LDWL[369],LDWL[368],LDWL[367],LDWL[366],LDWL[365],LDWL[364],LDWL[363],LDWL[362],LDWL[361],LDWL[360],LDWL[359],LDWL[358],LDWL[357],LDWL[356],LDWL[355],LDWL[354],LDWL[353],LDWL[352],LDWL[351],LDWL[350],LDWL[349],LDWL[348],LDWL[347],LDWL[346],LDWL[345],LDWL[344],LDWL[343],LDWL[342],LDWL[341],LDWL[340],LDWL[339],LDWL[338],LDWL[337],LDWL[336],LDWL[335],LDWL[334],LDWL[333],LDWL[332],LDWL[331],LDWL[330],LDWL[329],LDWL[328],LDWL[327],LDWL[326],LDWL[325],LDWL[324],LDWL[323],LDWL[322],LDWL[321],LDWL[320],LDWL[319],LDWL[318],LDWL[317],LDWL[316],LDWL[315],LDWL[314],LDWL[313],LDWL[312],LDWL[311],LDWL[310],LDWL[309],LDWL[308],LDWL[307],LDWL[306],LDWL[305],LDWL[304],LDWL[303],LDWL[302],LDWL[301],LDWL[300],LDWL[299],LDWL[298],LDWL[297],LDWL[296],LDWL[295],LDWL[294],LDWL[293],LDWL[292],LDWL[291],LDWL[290],LDWL[289],LDWL[288],LDWL[287],LDWL[286],LDWL[285],LDWL[284],LDWL[283],LDWL[282],LDWL[281],LDWL[280],LDWL[279],LDWL[278],LDWL[277],LDWL[276],LDWL[275],LDWL[274],LDWL[273],LDWL[272],LDWL[271],LDWL[270],LDWL[269],LDWL[268],LDWL[267],LDWL[266],LDWL[265],LDWL[264],LDWL[263],LDWL[262],LDWL[261],LDWL[260],LDWL[259],LDWL[258],LDWL[257],LDWL[256],LDWL[255],LDWL[254],LDWL[253],LDWL[252],LDWL[251],LDWL[250],LDWL[249],LDWL[248],LDWL[247],LDWL[246],LDWL[245],LDWL[244],LDWL[243],LDWL[242],LDWL[241],LDWL[240],LDWL[239],LDWL[238],LDWL[237],LDWL[236],LDWL[235],LDWL[234],LDWL[233],LDWL[232],LDWL[231],LDWL[230],LDWL[229],LDWL[228],LDWL[227],LDWL[226],LDWL[225],LDWL[224],LDWL[223],LDWL[222],LDWL[221],LDWL[220],LDWL[219],LDWL[218],LDWL[217],LDWL[216],LDWL[215],LDWL[214],LDWL[213],LDWL[212],LDWL[211],LDWL[210],LDWL[209],LDWL[208],LDWL[207],LDWL[206],LDWL[205],LDWL[204],LDWL[203],LDWL[202],LDWL[201],LDWL[200],LDWL[199],LDWL[198],LDWL[197],LDWL[196],LDWL[195],LDWL[194],LDWL[193],LDWL[192],LDWL[191],LDWL[190],LDWL[189],LDWL[188],LDWL[187],LDWL[186],LDWL[185],LDWL[184],LDWL[183],LDWL[182],LDWL[181],LDWL[180],LDWL[179],LDWL[178],LDWL[177],LDWL[176],LDWL[175],LDWL[174],LDWL[173],LDWL[172],LDWL[171],LDWL[170],LDWL[169],LDWL[168],LDWL[167],LDWL[166],LDWL[165],LDWL[164],LDWL[163],LDWL[162],LDWL[161],LDWL[160],LDWL[159],LDWL[158],LDWL[157],LDWL[156],LDWL[155],LDWL[154],LDWL[153],LDWL[152],LDWL[151],LDWL[150],LDWL[149],LDWL[148],LDWL[147],LDWL[146],LDWL[145],LDWL[144],LDWL[143],LDWL[142],LDWL[141],LDWL[140],LDWL[139],LDWL[138],LDWL[137],LDWL[136],LDWL[135],LDWL[134],LDWL[133],LDWL[132],LDWL[131],LDWL[130],LDWL[129],LDWL[128],LDWL[127],LDWL[126],LDWL[125],LDWL[124],LDWL[123],LDWL[122],LDWL[121],LDWL[120],LDWL[119],LDWL[118],LDWL[117],LDWL[116],LDWL[115],LDWL[114],LDWL[113],LDWL[112],LDWL[111],LDWL[110],LDWL[109],LDWL[108],LDWL[107],LDWL[106],LDWL[105],LDWL[104],LDWL[103],LDWL[102],LDWL[101],LDWL[100],LDWL[99],LDWL[98],LDWL[97],LDWL[96],LDWL[95],LDWL[94],LDWL[93],LDWL[92],LDWL[91],LDWL[90],LDWL[89],LDWL[88],LDWL[87],LDWL[86],LDWL[85],LDWL[84],LDWL[83],LDWL[82],LDWL[81],LDWL[80],LDWL[79],LDWL[78],LDWL[77],LDWL[76],LDWL[75],LDWL[74],LDWL[73],LDWL[72],LDWL[71],LDWL[70],LDWL[69],LDWL[68],LDWL[67],LDWL[66],LDWL[65],LDWL[64],LDWL[63],LDWL[62],LDWL[61],LDWL[60],LDWL[59],LDWL[58],LDWL[57],LDWL[56],LDWL[55],LDWL[54],LDWL[53],LDWL[52],LDWL[51],LDWL[50],LDWL[49],LDWL[48],LDWL[47],LDWL[46],LDWL[45],LDWL[44],LDWL[43],LDWL[42],LDWL[41],LDWL[40],LDWL[39],LDWL[38],LDWL[37],LDWL[36],LDWL[35],LDWL[34],LDWL[33],LDWL[32],LDWL[31],LDWL[30],LDWL[29],LDWL[28],LDWL[27],LDWL[26],LDWL[25],LDWL[24],LDWL[23],LDWL[22],LDWL[21],LDWL[20],LDWL[19],LDWL[18],LDWL[17],LDWL[16],LDWL[15],LDWL[14],LDWL[13],LDWL[12],LDWL[11],LDWL[10],LDWL[9],LDWL[8],LDWL[7],LDWL[6],LDWL[5],LDWL[4],LDWL[3],LDWL[2],LDWL[1],LDWL[0]
*.ipin vss
*.iopin LDBLREF
c1 LDBLREF 0 180f m=1
**** begin user architecture code
* PARASITICS


* reference bl


mr0 LDBLREF LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr1 LDBLREF LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr2 LDBLREF LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr3 LDBLREF LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr4 LDBLREF LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr5 LDBLREF LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr6 LDBLREF LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr7 LDBLREF LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr8 LDBLREF LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr9 LDBLREF LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
mr10 LDBLREF LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr11 LDBLREF LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr12 LDBLREF LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr13 LDBLREF LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr14 LDBLREF LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr15 LDBLREF LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr16 LDBLREF LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr17 LDBLREF LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr18 LDBLREF LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr19 LDBLREF LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr20 LDBLREF LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr21 LDBLREF LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr22 LDBLREF LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr23 LDBLREF LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr24 LDBLREF LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr25 LDBLREF LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr26 LDBLREF LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr27 LDBLREF LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr28 LDBLREF LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr29 LDBLREF LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr30 LDBLREF LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr31 LDBLREF LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr32 LDBLREF LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr33 LDBLREF LDWL[33] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr34 LDBLREF LDWL[34] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr35 LDBLREF LDWL[35] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr36 LDBLREF LDWL[36] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr37 LDBLREF LDWL[37] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr38 LDBLREF LDWL[38] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr39 LDBLREF LDWL[39] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr40 LDBLREF LDWL[40] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr41 LDBLREF LDWL[41] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr42 LDBLREF LDWL[42] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr43 LDBLREF LDWL[43] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr44 LDBLREF LDWL[44] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr45 LDBLREF LDWL[45] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr46 LDBLREF LDWL[46] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr47 LDBLREF LDWL[47] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr48 LDBLREF LDWL[48] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr49 LDBLREF LDWL[49] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr50 LDBLREF LDWL[50] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr51 LDBLREF LDWL[51] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr52 LDBLREF LDWL[52] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr53 LDBLREF LDWL[53] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr54 LDBLREF LDWL[54] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr55 LDBLREF LDWL[55] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr56 LDBLREF LDWL[56] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr57 LDBLREF LDWL[57] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr58 LDBLREF LDWL[58] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr59 LDBLREF LDWL[59] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr60 LDBLREF LDWL[60] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr61 LDBLREF LDWL[61] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr62 LDBLREF LDWL[62] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr63 LDBLREF LDWL[63] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr64 LDBLREF LDWL[64] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr65 LDBLREF LDWL[65] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr66 LDBLREF LDWL[66] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr67 LDBLREF LDWL[67] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr68 LDBLREF LDWL[68] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr69 LDBLREF LDWL[69] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr70 LDBLREF LDWL[70] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr71 LDBLREF LDWL[71] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr72 LDBLREF LDWL[72] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr73 LDBLREF LDWL[73] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr74 LDBLREF LDWL[74] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr75 LDBLREF LDWL[75] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr76 LDBLREF LDWL[76] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr77 LDBLREF LDWL[77] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr78 LDBLREF LDWL[78] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr79 LDBLREF LDWL[79] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr80 LDBLREF LDWL[80] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr81 LDBLREF LDWL[81] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr82 LDBLREF LDWL[82] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr83 LDBLREF LDWL[83] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr84 LDBLREF LDWL[84] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr85 LDBLREF LDWL[85] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr86 LDBLREF LDWL[86] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr87 LDBLREF LDWL[87] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr88 LDBLREF LDWL[88] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr89 LDBLREF LDWL[89] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr90 LDBLREF LDWL[90] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr91 LDBLREF LDWL[91] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr92 LDBLREF LDWL[92] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr93 LDBLREF LDWL[93] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr94 LDBLREF LDWL[94] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr95 LDBLREF LDWL[95] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr96 LDBLREF LDWL[96] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr97 LDBLREF LDWL[97] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr98 LDBLREF LDWL[98] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr99 LDBLREF LDWL[99] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr100 LDBLREF LDWL[100] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr101 LDBLREF LDWL[101] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr102 LDBLREF LDWL[102] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr103 LDBLREF LDWL[103] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr104 LDBLREF LDWL[104] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr105 LDBLREF LDWL[105] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr106 LDBLREF LDWL[106] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr107 LDBLREF LDWL[107] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr108 LDBLREF LDWL[108] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr109 LDBLREF LDWL[109] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr110 LDBLREF LDWL[110] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr111 LDBLREF LDWL[111] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr112 LDBLREF LDWL[112] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr113 LDBLREF LDWL[113] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr114 LDBLREF LDWL[114] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr115 LDBLREF LDWL[115] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr116 LDBLREF LDWL[116] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr117 LDBLREF LDWL[117] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr118 LDBLREF LDWL[118] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr119 LDBLREF LDWL[119] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr120 LDBLREF LDWL[120] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr121 LDBLREF LDWL[121] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr122 LDBLREF LDWL[122] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr123 LDBLREF LDWL[123] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr124 LDBLREF LDWL[124] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr125 LDBLREF LDWL[125] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr126 LDBLREF LDWL[126] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr127 LDBLREF LDWL[127] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr128 LDBLREF LDWL[128] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr129 LDBLREF LDWL[129] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr130 LDBLREF LDWL[130] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr131 LDBLREF LDWL[131] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr132 LDBLREF LDWL[132] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr133 LDBLREF LDWL[133] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr134 LDBLREF LDWL[134] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr135 LDBLREF LDWL[135] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr136 LDBLREF LDWL[136] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr137 LDBLREF LDWL[137] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr138 LDBLREF LDWL[138] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr139 LDBLREF LDWL[139] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr140 LDBLREF LDWL[140] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr141 LDBLREF LDWL[141] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr142 LDBLREF LDWL[142] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr143 LDBLREF LDWL[143] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr144 LDBLREF LDWL[144] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr145 LDBLREF LDWL[145] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr146 LDBLREF LDWL[146] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr147 LDBLREF LDWL[147] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr148 LDBLREF LDWL[148] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr149 LDBLREF LDWL[149] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr150 LDBLREF LDWL[150] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr151 LDBLREF LDWL[151] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr152 LDBLREF LDWL[152] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr153 LDBLREF LDWL[153] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr154 LDBLREF LDWL[154] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr155 LDBLREF LDWL[155] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr156 LDBLREF LDWL[156] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr157 LDBLREF LDWL[157] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr158 LDBLREF LDWL[158] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr159 LDBLREF LDWL[159] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr160 LDBLREF LDWL[160] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr161 LDBLREF LDWL[161] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr162 LDBLREF LDWL[162] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr163 LDBLREF LDWL[163] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr164 LDBLREF LDWL[164] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr165 LDBLREF LDWL[165] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr166 LDBLREF LDWL[166] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr167 LDBLREF LDWL[167] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr168 LDBLREF LDWL[168] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr169 LDBLREF LDWL[169] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr170 LDBLREF LDWL[170] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr171 LDBLREF LDWL[171] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr172 LDBLREF LDWL[172] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr173 LDBLREF LDWL[173] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr174 LDBLREF LDWL[174] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr175 LDBLREF LDWL[175] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr176 LDBLREF LDWL[176] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr177 LDBLREF LDWL[177] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr178 LDBLREF LDWL[178] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr179 LDBLREF LDWL[179] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr180 LDBLREF LDWL[180] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr181 LDBLREF LDWL[181] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr182 LDBLREF LDWL[182] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr183 LDBLREF LDWL[183] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr184 LDBLREF LDWL[184] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr185 LDBLREF LDWL[185] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr186 LDBLREF LDWL[186] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr187 LDBLREF LDWL[187] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr188 LDBLREF LDWL[188] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr189 LDBLREF LDWL[189] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr190 LDBLREF LDWL[190] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr191 LDBLREF LDWL[191] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr192 LDBLREF LDWL[192] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr193 LDBLREF LDWL[193] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr194 LDBLREF LDWL[194] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr195 LDBLREF LDWL[195] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr196 LDBLREF LDWL[196] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr197 LDBLREF LDWL[197] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr198 LDBLREF LDWL[198] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr199 LDBLREF LDWL[199] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr200 LDBLREF LDWL[200] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr201 LDBLREF LDWL[201] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr202 LDBLREF LDWL[202] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr203 LDBLREF LDWL[203] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr204 LDBLREF LDWL[204] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr205 LDBLREF LDWL[205] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr206 LDBLREF LDWL[206] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr207 LDBLREF LDWL[207] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr208 LDBLREF LDWL[208] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr209 LDBLREF LDWL[209] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr210 LDBLREF LDWL[210] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr211 LDBLREF LDWL[211] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr212 LDBLREF LDWL[212] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr213 LDBLREF LDWL[213] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr214 LDBLREF LDWL[214] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr215 LDBLREF LDWL[215] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr216 LDBLREF LDWL[216] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr217 LDBLREF LDWL[217] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr218 LDBLREF LDWL[218] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr219 LDBLREF LDWL[219] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr220 LDBLREF LDWL[220] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr221 LDBLREF LDWL[221] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr222 LDBLREF LDWL[222] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr223 LDBLREF LDWL[223] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr224 LDBLREF LDWL[224] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr225 LDBLREF LDWL[225] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr226 LDBLREF LDWL[226] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr227 LDBLREF LDWL[227] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr228 LDBLREF LDWL[228] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr229 LDBLREF LDWL[229] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr230 LDBLREF LDWL[230] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr231 LDBLREF LDWL[231] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr232 LDBLREF LDWL[232] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr233 LDBLREF LDWL[233] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr234 LDBLREF LDWL[234] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr235 LDBLREF LDWL[235] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr236 LDBLREF LDWL[236] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr237 LDBLREF LDWL[237] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr238 LDBLREF LDWL[238] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr239 LDBLREF LDWL[239] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr240 LDBLREF LDWL[240] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr241 LDBLREF LDWL[241] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr242 LDBLREF LDWL[242] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr243 LDBLREF LDWL[243] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr244 LDBLREF LDWL[244] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr245 LDBLREF LDWL[245] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr246 LDBLREF LDWL[246] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr247 LDBLREF LDWL[247] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr248 LDBLREF LDWL[248] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr249 LDBLREF LDWL[249] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr250 LDBLREF LDWL[250] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr251 LDBLREF LDWL[251] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr252 LDBLREF LDWL[252] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr253 LDBLREF LDWL[253] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr254 LDBLREF LDWL[254] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr255 LDBLREF LDWL[255] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr256 LDBLREF LDWL[256] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr257 LDBLREF LDWL[257] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr258 LDBLREF LDWL[258] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr259 LDBLREF LDWL[259] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr260 LDBLREF LDWL[260] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr261 LDBLREF LDWL[261] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr262 LDBLREF LDWL[262] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr263 LDBLREF LDWL[263] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr264 LDBLREF LDWL[264] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr265 LDBLREF LDWL[265] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr266 LDBLREF LDWL[266] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr267 LDBLREF LDWL[267] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr268 LDBLREF LDWL[268] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr269 LDBLREF LDWL[269] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr270 LDBLREF LDWL[270] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr271 LDBLREF LDWL[271] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr272 LDBLREF LDWL[272] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr273 LDBLREF LDWL[273] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr274 LDBLREF LDWL[274] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr275 LDBLREF LDWL[275] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr276 LDBLREF LDWL[276] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr277 LDBLREF LDWL[277] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr278 LDBLREF LDWL[278] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr279 LDBLREF LDWL[279] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr280 LDBLREF LDWL[280] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr281 LDBLREF LDWL[281] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr282 LDBLREF LDWL[282] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr283 LDBLREF LDWL[283] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr284 LDBLREF LDWL[284] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr285 LDBLREF LDWL[285] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr286 LDBLREF LDWL[286] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr287 LDBLREF LDWL[287] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr288 LDBLREF LDWL[288] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr289 LDBLREF LDWL[289] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr290 LDBLREF LDWL[290] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr291 LDBLREF LDWL[291] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr292 LDBLREF LDWL[292] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr293 LDBLREF LDWL[293] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr294 LDBLREF LDWL[294] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr295 LDBLREF LDWL[295] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr296 LDBLREF LDWL[296] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr297 LDBLREF LDWL[297] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr298 LDBLREF LDWL[298] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr299 LDBLREF LDWL[299] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr300 LDBLREF LDWL[300] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr301 LDBLREF LDWL[301] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr302 LDBLREF LDWL[302] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr303 LDBLREF LDWL[303] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr304 LDBLREF LDWL[304] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr305 LDBLREF LDWL[305] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr306 LDBLREF LDWL[306] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr307 LDBLREF LDWL[307] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr308 LDBLREF LDWL[308] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr309 LDBLREF LDWL[309] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr310 LDBLREF LDWL[310] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr311 LDBLREF LDWL[311] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr312 LDBLREF LDWL[312] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr313 LDBLREF LDWL[313] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr314 LDBLREF LDWL[314] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr315 LDBLREF LDWL[315] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr316 LDBLREF LDWL[316] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr317 LDBLREF LDWL[317] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr318 LDBLREF LDWL[318] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr319 LDBLREF LDWL[319] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr320 LDBLREF LDWL[320] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr321 LDBLREF LDWL[321] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr322 LDBLREF LDWL[322] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr323 LDBLREF LDWL[323] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr324 LDBLREF LDWL[324] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr325 LDBLREF LDWL[325] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr326 LDBLREF LDWL[326] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr327 LDBLREF LDWL[327] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr328 LDBLREF LDWL[328] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr329 LDBLREF LDWL[329] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr330 LDBLREF LDWL[330] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr331 LDBLREF LDWL[331] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr332 LDBLREF LDWL[332] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr333 LDBLREF LDWL[333] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr334 LDBLREF LDWL[334] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr335 LDBLREF LDWL[335] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr336 LDBLREF LDWL[336] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr337 LDBLREF LDWL[337] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr338 LDBLREF LDWL[338] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr339 LDBLREF LDWL[339] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr340 LDBLREF LDWL[340] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr341 LDBLREF LDWL[341] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr342 LDBLREF LDWL[342] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr343 LDBLREF LDWL[343] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr344 LDBLREF LDWL[344] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr345 LDBLREF LDWL[345] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr346 LDBLREF LDWL[346] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr347 LDBLREF LDWL[347] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr348 LDBLREF LDWL[348] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr349 LDBLREF LDWL[349] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr350 LDBLREF LDWL[350] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr351 LDBLREF LDWL[351] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr352 LDBLREF LDWL[352] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr353 LDBLREF LDWL[353] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr354 LDBLREF LDWL[354] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr355 LDBLREF LDWL[355] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr356 LDBLREF LDWL[356] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr357 LDBLREF LDWL[357] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr358 LDBLREF LDWL[358] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr359 LDBLREF LDWL[359] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr360 LDBLREF LDWL[360] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr361 LDBLREF LDWL[361] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr362 LDBLREF LDWL[362] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr363 LDBLREF LDWL[363] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr364 LDBLREF LDWL[364] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr365 LDBLREF LDWL[365] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr366 LDBLREF LDWL[366] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr367 LDBLREF LDWL[367] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr368 LDBLREF LDWL[368] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr369 LDBLREF LDWL[369] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr370 LDBLREF LDWL[370] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr371 LDBLREF LDWL[371] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr372 LDBLREF LDWL[372] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr373 LDBLREF LDWL[373] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr374 LDBLREF LDWL[374] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr375 LDBLREF LDWL[375] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr376 LDBLREF LDWL[376] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr377 LDBLREF LDWL[377] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr378 LDBLREF LDWL[378] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr379 LDBLREF LDWL[379] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr380 LDBLREF LDWL[380] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr381 LDBLREF LDWL[381] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr382 LDBLREF LDWL[382] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr383 LDBLREF LDWL[383] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr384 LDBLREF LDWL[384] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr385 LDBLREF LDWL[385] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr386 LDBLREF LDWL[386] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr387 LDBLREF LDWL[387] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr388 LDBLREF LDWL[388] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr389 LDBLREF LDWL[389] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr390 LDBLREF LDWL[390] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr391 LDBLREF LDWL[391] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr392 LDBLREF LDWL[392] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr393 LDBLREF LDWL[393] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr394 LDBLREF LDWL[394] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr395 LDBLREF LDWL[395] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr396 LDBLREF LDWL[396] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr397 LDBLREF LDWL[397] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr398 LDBLREF LDWL[398] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr399 LDBLREF LDWL[399] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr400 LDBLREF LDWL[400] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr401 LDBLREF LDWL[401] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr402 LDBLREF LDWL[402] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr403 LDBLREF LDWL[403] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr404 LDBLREF LDWL[404] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr405 LDBLREF LDWL[405] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr406 LDBLREF LDWL[406] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr407 LDBLREF LDWL[407] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr408 LDBLREF LDWL[408] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr409 LDBLREF LDWL[409] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr410 LDBLREF LDWL[410] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr411 LDBLREF LDWL[411] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr412 LDBLREF LDWL[412] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr413 LDBLREF LDWL[413] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr414 LDBLREF LDWL[414] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr415 LDBLREF LDWL[415] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr416 LDBLREF LDWL[416] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr417 LDBLREF LDWL[417] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr418 LDBLREF LDWL[418] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr419 LDBLREF LDWL[419] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr420 LDBLREF LDWL[420] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr421 LDBLREF LDWL[421] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr422 LDBLREF LDWL[422] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr423 LDBLREF LDWL[423] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr424 LDBLREF LDWL[424] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr425 LDBLREF LDWL[425] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr426 LDBLREF LDWL[426] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr427 LDBLREF LDWL[427] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr428 LDBLREF LDWL[428] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr429 LDBLREF LDWL[429] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr430 LDBLREF LDWL[430] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr431 LDBLREF LDWL[431] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr432 LDBLREF LDWL[432] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr433 LDBLREF LDWL[433] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr434 LDBLREF LDWL[434] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr435 LDBLREF LDWL[435] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr436 LDBLREF LDWL[436] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr437 LDBLREF LDWL[437] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr438 LDBLREF LDWL[438] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr439 LDBLREF LDWL[439] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr440 LDBLREF LDWL[440] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr441 LDBLREF LDWL[441] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr442 LDBLREF LDWL[442] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr443 LDBLREF LDWL[443] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr444 LDBLREF LDWL[444] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr445 LDBLREF LDWL[445] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr446 LDBLREF LDWL[446] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr447 LDBLREF LDWL[447] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr448 LDBLREF LDWL[448] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr449 LDBLREF LDWL[449] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr450 LDBLREF LDWL[450] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr451 LDBLREF LDWL[451] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr452 LDBLREF LDWL[452] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr453 LDBLREF LDWL[453] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr454 LDBLREF LDWL[454] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr455 LDBLREF LDWL[455] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr456 LDBLREF LDWL[456] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr457 LDBLREF LDWL[457] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr458 LDBLREF LDWL[458] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr459 LDBLREF LDWL[459] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr460 LDBLREF LDWL[460] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr461 LDBLREF LDWL[461] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr462 LDBLREF LDWL[462] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr463 LDBLREF LDWL[463] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr464 LDBLREF LDWL[464] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr465 LDBLREF LDWL[465] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr466 LDBLREF LDWL[466] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr467 LDBLREF LDWL[467] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr468 LDBLREF LDWL[468] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr469 LDBLREF LDWL[469] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr470 LDBLREF LDWL[470] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr471 LDBLREF LDWL[471] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr472 LDBLREF LDWL[472] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr473 LDBLREF LDWL[473] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr474 LDBLREF LDWL[474] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr475 LDBLREF LDWL[475] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr476 LDBLREF LDWL[476] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr477 LDBLREF LDWL[477] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr478 LDBLREF LDWL[478] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr479 LDBLREF LDWL[479] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr480 LDBLREF LDWL[480] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr481 LDBLREF LDWL[481] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr482 LDBLREF LDWL[482] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr483 LDBLREF LDWL[483] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr484 LDBLREF LDWL[484] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr485 LDBLREF LDWL[485] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr486 LDBLREF LDWL[486] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr487 LDBLREF LDWL[487] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr488 LDBLREF LDWL[488] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr489 LDBLREF LDWL[489] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr490 LDBLREF LDWL[490] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr491 LDBLREF LDWL[491] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr492 LDBLREF LDWL[492] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr493 LDBLREF LDWL[493] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr494 LDBLREF LDWL[494] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr495 LDBLREF LDWL[495] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr496 LDBLREF LDWL[496] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr497 LDBLREF LDWL[497] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr498 LDBLREF LDWL[498] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr499 LDBLREF LDWL[499] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr500 LDBLREF LDWL[500] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr501 LDBLREF LDWL[501] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr502 LDBLREF LDWL[502] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr503 LDBLREF LDWL[503] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr504 LDBLREF LDWL[504] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr505 LDBLREF LDWL[505] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr506 LDBLREF LDWL[506] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr507 LDBLREF LDWL[507] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr508 LDBLREF LDWL[508] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr509 LDBLREF LDWL[509] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr510 LDBLREF LDWL[510] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
mr511 LDBLREF LDWL[511] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1

* /reference bl

* last bitline


ml0 VSS LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml1 VSS LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml2 VSS LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml3 VSS LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml4 VSS LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml5 VSS LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml6 VSS LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml7 VSS LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml8 VSS LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml9 VSS LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml10 VSS LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml11 VSS LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml12 VSS LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml13 VSS LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml14 VSS LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml15 VSS LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml16 VSS LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml17 VSS LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml18 VSS LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml19 VSS LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml20 VSS LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml21 VSS LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml22 VSS LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml23 VSS LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml24 VSS LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml25 VSS LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml26 VSS LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml27 VSS LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml28 VSS LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml29 VSS LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml30 VSS LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml31 VSS LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml32 VSS LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml33 VSS LDWL[33] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml34 VSS LDWL[34] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml35 VSS LDWL[35] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml36 VSS LDWL[36] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml37 VSS LDWL[37] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml38 VSS LDWL[38] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml39 VSS LDWL[39] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml40 VSS LDWL[40] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml41 VSS LDWL[41] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml42 VSS LDWL[42] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml43 VSS LDWL[43] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml44 VSS LDWL[44] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml45 VSS LDWL[45] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml46 VSS LDWL[46] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml47 VSS LDWL[47] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml48 VSS LDWL[48] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml49 VSS LDWL[49] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml50 VSS LDWL[50] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml51 VSS LDWL[51] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml52 VSS LDWL[52] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml53 VSS LDWL[53] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml54 VSS LDWL[54] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml55 VSS LDWL[55] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml56 VSS LDWL[56] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml57 VSS LDWL[57] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml58 VSS LDWL[58] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml59 VSS LDWL[59] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml60 VSS LDWL[60] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml61 VSS LDWL[61] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml62 VSS LDWL[62] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml63 VSS LDWL[63] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml64 VSS LDWL[64] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml65 VSS LDWL[65] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml66 VSS LDWL[66] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml67 VSS LDWL[67] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml68 VSS LDWL[68] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml69 VSS LDWL[69] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml70 VSS LDWL[70] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml71 VSS LDWL[71] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml72 VSS LDWL[72] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml73 VSS LDWL[73] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml74 VSS LDWL[74] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml75 VSS LDWL[75] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml76 VSS LDWL[76] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml77 VSS LDWL[77] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml78 VSS LDWL[78] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml79 VSS LDWL[79] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml80 VSS LDWL[80] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml81 VSS LDWL[81] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml82 VSS LDWL[82] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml83 VSS LDWL[83] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml84 VSS LDWL[84] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml85 VSS LDWL[85] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml86 VSS LDWL[86] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml87 VSS LDWL[87] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml88 VSS LDWL[88] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml89 VSS LDWL[89] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml90 VSS LDWL[90] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml91 VSS LDWL[91] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml92 VSS LDWL[92] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml93 VSS LDWL[93] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml94 VSS LDWL[94] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml95 VSS LDWL[95] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml96 VSS LDWL[96] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml97 VSS LDWL[97] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml98 VSS LDWL[98] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml99 VSS LDWL[99] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml100 VSS LDWL[100] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml101 VSS LDWL[101] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml102 VSS LDWL[102] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml103 VSS LDWL[103] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml104 VSS LDWL[104] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml105 VSS LDWL[105] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml106 VSS LDWL[106] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml107 VSS LDWL[107] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml108 VSS LDWL[108] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml109 VSS LDWL[109] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml110 VSS LDWL[110] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml111 VSS LDWL[111] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml112 VSS LDWL[112] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml113 VSS LDWL[113] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml114 VSS LDWL[114] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml115 VSS LDWL[115] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml116 VSS LDWL[116] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml117 VSS LDWL[117] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml118 VSS LDWL[118] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml119 VSS LDWL[119] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml120 VSS LDWL[120] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml121 VSS LDWL[121] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml122 VSS LDWL[122] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml123 VSS LDWL[123] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml124 VSS LDWL[124] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml125 VSS LDWL[125] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml126 VSS LDWL[126] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml127 VSS LDWL[127] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml128 VSS LDWL[128] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml129 VSS LDWL[129] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml130 VSS LDWL[130] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml131 VSS LDWL[131] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml132 VSS LDWL[132] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml133 VSS LDWL[133] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml134 VSS LDWL[134] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml135 VSS LDWL[135] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml136 VSS LDWL[136] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml137 VSS LDWL[137] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml138 VSS LDWL[138] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml139 VSS LDWL[139] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml140 VSS LDWL[140] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml141 VSS LDWL[141] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml142 VSS LDWL[142] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml143 VSS LDWL[143] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml144 VSS LDWL[144] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml145 VSS LDWL[145] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml146 VSS LDWL[146] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml147 VSS LDWL[147] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml148 VSS LDWL[148] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml149 VSS LDWL[149] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml150 VSS LDWL[150] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml151 VSS LDWL[151] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml152 VSS LDWL[152] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml153 VSS LDWL[153] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml154 VSS LDWL[154] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml155 VSS LDWL[155] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml156 VSS LDWL[156] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml157 VSS LDWL[157] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml158 VSS LDWL[158] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml159 VSS LDWL[159] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml160 VSS LDWL[160] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml161 VSS LDWL[161] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml162 VSS LDWL[162] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml163 VSS LDWL[163] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml164 VSS LDWL[164] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml165 VSS LDWL[165] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml166 VSS LDWL[166] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml167 VSS LDWL[167] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml168 VSS LDWL[168] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml169 VSS LDWL[169] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml170 VSS LDWL[170] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml171 VSS LDWL[171] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml172 VSS LDWL[172] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml173 VSS LDWL[173] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml174 VSS LDWL[174] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml175 VSS LDWL[175] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml176 VSS LDWL[176] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml177 VSS LDWL[177] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml178 VSS LDWL[178] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml179 VSS LDWL[179] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml180 VSS LDWL[180] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml181 VSS LDWL[181] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml182 VSS LDWL[182] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml183 VSS LDWL[183] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml184 VSS LDWL[184] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml185 VSS LDWL[185] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml186 VSS LDWL[186] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml187 VSS LDWL[187] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml188 VSS LDWL[188] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml189 VSS LDWL[189] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml190 VSS LDWL[190] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml191 VSS LDWL[191] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml192 VSS LDWL[192] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml193 VSS LDWL[193] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml194 VSS LDWL[194] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml195 VSS LDWL[195] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml196 VSS LDWL[196] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml197 VSS LDWL[197] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml198 VSS LDWL[198] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml199 VSS LDWL[199] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml200 VSS LDWL[200] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml201 VSS LDWL[201] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml202 VSS LDWL[202] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml203 VSS LDWL[203] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml204 VSS LDWL[204] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml205 VSS LDWL[205] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml206 VSS LDWL[206] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml207 VSS LDWL[207] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml208 VSS LDWL[208] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml209 VSS LDWL[209] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml210 VSS LDWL[210] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml211 VSS LDWL[211] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml212 VSS LDWL[212] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml213 VSS LDWL[213] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml214 VSS LDWL[214] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml215 VSS LDWL[215] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml216 VSS LDWL[216] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml217 VSS LDWL[217] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml218 VSS LDWL[218] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml219 VSS LDWL[219] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml220 VSS LDWL[220] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml221 VSS LDWL[221] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml222 VSS LDWL[222] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml223 VSS LDWL[223] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml224 VSS LDWL[224] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml225 VSS LDWL[225] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml226 VSS LDWL[226] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml227 VSS LDWL[227] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml228 VSS LDWL[228] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml229 VSS LDWL[229] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml230 VSS LDWL[230] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml231 VSS LDWL[231] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml232 VSS LDWL[232] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml233 VSS LDWL[233] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml234 VSS LDWL[234] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml235 VSS LDWL[235] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml236 VSS LDWL[236] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml237 VSS LDWL[237] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml238 VSS LDWL[238] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml239 VSS LDWL[239] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml240 VSS LDWL[240] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml241 VSS LDWL[241] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml242 VSS LDWL[242] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml243 VSS LDWL[243] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml244 VSS LDWL[244] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml245 VSS LDWL[245] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml246 VSS LDWL[246] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml247 VSS LDWL[247] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml248 VSS LDWL[248] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml249 VSS LDWL[249] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml250 VSS LDWL[250] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml251 VSS LDWL[251] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml252 VSS LDWL[252] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml253 VSS LDWL[253] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml254 VSS LDWL[254] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml255 VSS LDWL[255] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml256 VSS LDWL[256] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml257 VSS LDWL[257] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml258 VSS LDWL[258] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml259 VSS LDWL[259] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml260 VSS LDWL[260] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml261 VSS LDWL[261] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml262 VSS LDWL[262] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml263 VSS LDWL[263] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml264 VSS LDWL[264] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml265 VSS LDWL[265] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml266 VSS LDWL[266] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml267 VSS LDWL[267] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml268 VSS LDWL[268] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml269 VSS LDWL[269] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml270 VSS LDWL[270] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml271 VSS LDWL[271] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml272 VSS LDWL[272] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml273 VSS LDWL[273] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml274 VSS LDWL[274] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml275 VSS LDWL[275] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml276 VSS LDWL[276] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml277 VSS LDWL[277] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml278 VSS LDWL[278] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml279 VSS LDWL[279] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml280 VSS LDWL[280] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml281 VSS LDWL[281] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml282 VSS LDWL[282] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml283 VSS LDWL[283] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml284 VSS LDWL[284] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml285 VSS LDWL[285] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml286 VSS LDWL[286] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml287 VSS LDWL[287] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml288 VSS LDWL[288] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml289 VSS LDWL[289] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml290 VSS LDWL[290] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml291 VSS LDWL[291] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml292 VSS LDWL[292] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml293 VSS LDWL[293] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml294 VSS LDWL[294] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml295 VSS LDWL[295] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml296 VSS LDWL[296] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml297 VSS LDWL[297] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml298 VSS LDWL[298] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml299 VSS LDWL[299] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml300 VSS LDWL[300] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml301 VSS LDWL[301] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml302 VSS LDWL[302] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml303 VSS LDWL[303] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml304 VSS LDWL[304] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml305 VSS LDWL[305] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml306 VSS LDWL[306] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml307 VSS LDWL[307] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml308 VSS LDWL[308] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml309 VSS LDWL[309] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml310 VSS LDWL[310] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml311 VSS LDWL[311] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml312 VSS LDWL[312] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml313 VSS LDWL[313] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml314 VSS LDWL[314] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml315 VSS LDWL[315] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml316 VSS LDWL[316] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml317 VSS LDWL[317] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml318 VSS LDWL[318] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml319 VSS LDWL[319] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml320 VSS LDWL[320] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml321 VSS LDWL[321] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml322 VSS LDWL[322] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml323 VSS LDWL[323] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml324 VSS LDWL[324] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml325 VSS LDWL[325] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml326 VSS LDWL[326] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml327 VSS LDWL[327] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml328 VSS LDWL[328] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml329 VSS LDWL[329] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml330 VSS LDWL[330] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml331 VSS LDWL[331] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml332 VSS LDWL[332] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml333 VSS LDWL[333] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml334 VSS LDWL[334] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml335 VSS LDWL[335] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml336 VSS LDWL[336] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml337 VSS LDWL[337] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml338 VSS LDWL[338] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml339 VSS LDWL[339] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml340 VSS LDWL[340] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml341 VSS LDWL[341] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml342 VSS LDWL[342] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml343 VSS LDWL[343] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml344 VSS LDWL[344] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml345 VSS LDWL[345] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml346 VSS LDWL[346] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml347 VSS LDWL[347] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml348 VSS LDWL[348] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml349 VSS LDWL[349] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml350 VSS LDWL[350] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml351 VSS LDWL[351] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml352 VSS LDWL[352] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml353 VSS LDWL[353] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml354 VSS LDWL[354] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml355 VSS LDWL[355] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml356 VSS LDWL[356] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml357 VSS LDWL[357] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml358 VSS LDWL[358] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml359 VSS LDWL[359] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml360 VSS LDWL[360] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml361 VSS LDWL[361] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml362 VSS LDWL[362] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml363 VSS LDWL[363] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml364 VSS LDWL[364] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml365 VSS LDWL[365] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml366 VSS LDWL[366] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml367 VSS LDWL[367] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml368 VSS LDWL[368] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml369 VSS LDWL[369] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml370 VSS LDWL[370] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml371 VSS LDWL[371] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml372 VSS LDWL[372] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml373 VSS LDWL[373] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml374 VSS LDWL[374] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml375 VSS LDWL[375] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml376 VSS LDWL[376] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml377 VSS LDWL[377] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml378 VSS LDWL[378] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml379 VSS LDWL[379] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml380 VSS LDWL[380] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml381 VSS LDWL[381] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml382 VSS LDWL[382] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml383 VSS LDWL[383] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml384 VSS LDWL[384] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml385 VSS LDWL[385] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml386 VSS LDWL[386] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml387 VSS LDWL[387] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml388 VSS LDWL[388] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml389 VSS LDWL[389] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml390 VSS LDWL[390] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml391 VSS LDWL[391] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml392 VSS LDWL[392] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml393 VSS LDWL[393] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml394 VSS LDWL[394] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml395 VSS LDWL[395] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml396 VSS LDWL[396] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml397 VSS LDWL[397] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml398 VSS LDWL[398] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml399 VSS LDWL[399] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml400 VSS LDWL[400] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml401 VSS LDWL[401] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml402 VSS LDWL[402] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml403 VSS LDWL[403] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml404 VSS LDWL[404] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml405 VSS LDWL[405] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml406 VSS LDWL[406] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml407 VSS LDWL[407] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml408 VSS LDWL[408] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml409 VSS LDWL[409] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml410 VSS LDWL[410] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml411 VSS LDWL[411] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml412 VSS LDWL[412] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml413 VSS LDWL[413] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml414 VSS LDWL[414] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml415 VSS LDWL[415] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml416 VSS LDWL[416] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml417 VSS LDWL[417] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml418 VSS LDWL[418] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml419 VSS LDWL[419] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml420 VSS LDWL[420] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml421 VSS LDWL[421] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml422 VSS LDWL[422] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml423 VSS LDWL[423] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml424 VSS LDWL[424] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml425 VSS LDWL[425] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml426 VSS LDWL[426] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml427 VSS LDWL[427] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml428 VSS LDWL[428] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml429 VSS LDWL[429] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml430 VSS LDWL[430] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml431 VSS LDWL[431] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml432 VSS LDWL[432] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml433 VSS LDWL[433] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml434 VSS LDWL[434] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml435 VSS LDWL[435] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml436 VSS LDWL[436] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml437 VSS LDWL[437] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml438 VSS LDWL[438] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml439 VSS LDWL[439] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml440 VSS LDWL[440] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml441 VSS LDWL[441] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml442 VSS LDWL[442] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml443 VSS LDWL[443] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml444 VSS LDWL[444] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml445 VSS LDWL[445] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml446 VSS LDWL[446] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml447 VSS LDWL[447] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml448 VSS LDWL[448] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml449 VSS LDWL[449] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml450 VSS LDWL[450] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml451 VSS LDWL[451] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml452 VSS LDWL[452] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml453 VSS LDWL[453] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml454 VSS LDWL[454] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml455 VSS LDWL[455] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml456 VSS LDWL[456] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml457 VSS LDWL[457] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml458 VSS LDWL[458] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml459 VSS LDWL[459] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml460 VSS LDWL[460] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml461 VSS LDWL[461] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml462 VSS LDWL[462] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml463 VSS LDWL[463] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml464 VSS LDWL[464] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml465 VSS LDWL[465] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml466 VSS LDWL[466] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml467 VSS LDWL[467] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml468 VSS LDWL[468] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml469 VSS LDWL[469] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml470 VSS LDWL[470] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml471 VSS LDWL[471] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml472 VSS LDWL[472] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml473 VSS LDWL[473] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml474 VSS LDWL[474] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml475 VSS LDWL[475] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml476 VSS LDWL[476] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml477 VSS LDWL[477] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml478 VSS LDWL[478] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml479 VSS LDWL[479] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml480 VSS LDWL[480] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml481 VSS LDWL[481] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml482 VSS LDWL[482] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml483 VSS LDWL[483] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml484 VSS LDWL[484] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml485 VSS LDWL[485] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml486 VSS LDWL[486] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml487 VSS LDWL[487] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml488 VSS LDWL[488] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml489 VSS LDWL[489] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml490 VSS LDWL[490] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml491 VSS LDWL[491] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml492 VSS LDWL[492] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml493 VSS LDWL[493] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml494 VSS LDWL[494] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml495 VSS LDWL[495] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml496 VSS LDWL[496] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml497 VSS LDWL[497] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml498 VSS LDWL[498] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml499 VSS LDWL[499] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml500 VSS LDWL[500] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml501 VSS LDWL[501] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml502 VSS LDWL[502] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml503 VSS LDWL[503] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml504 VSS LDWL[504] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml505 VSS LDWL[505] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml506 VSS LDWL[506] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml507 VSS LDWL[507] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml508 VSS LDWL[508] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml509 VSS LDWL[509] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml510 VSS LDWL[510] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
ml511 VSS LDWL[511] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1

* /last bitline



**** end user architecture code
.ends


* expanding   symbol:  rom2_col_prech.sym # of pins=3
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_col_prech.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_col_prech.sch
.subckt rom2_col_prech  LDPRECH LDBL vss
*.iopin LDBL
*.ipin LDPRECH
*.ipin vss
m0 vss LDPRECH LDBL 0 cmosn w=6u l=2.4u ad='6u *4.4u' as='6u *4.4u' pd='6u *2 + 8.8u' ps='6u *2 + 8.8u'
+ m=1
.ends


* expanding   symbol:  rom3_array.sym # of pins=3
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom3_array.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom3_array.sch
.subckt rom3_array  LDWL[511] LDWL[510] LDWL[509] LDWL[508] LDWL[507] LDWL[506] LDWL[505] LDWL[504]
+ LDWL[503] LDWL[502] LDWL[501] LDWL[500] LDWL[499] LDWL[498] LDWL[497] LDWL[496] LDWL[495] LDWL[494] LDWL[493]
+ LDWL[492] LDWL[491] LDWL[490] LDWL[489] LDWL[488] LDWL[487] LDWL[486] LDWL[485] LDWL[484] LDWL[483] LDWL[482]
+ LDWL[481] LDWL[480] LDWL[479] LDWL[478] LDWL[477] LDWL[476] LDWL[475] LDWL[474] LDWL[473] LDWL[472] LDWL[471]
+ LDWL[470] LDWL[469] LDWL[468] LDWL[467] LDWL[466] LDWL[465] LDWL[464] LDWL[463] LDWL[462] LDWL[461] LDWL[460]
+ LDWL[459] LDWL[458] LDWL[457] LDWL[456] LDWL[455] LDWL[454] LDWL[453] LDWL[452] LDWL[451] LDWL[450] LDWL[449]
+ LDWL[448] LDWL[447] LDWL[446] LDWL[445] LDWL[444] LDWL[443] LDWL[442] LDWL[441] LDWL[440] LDWL[439] LDWL[438]
+ LDWL[437] LDWL[436] LDWL[435] LDWL[434] LDWL[433] LDWL[432] LDWL[431] LDWL[430] LDWL[429] LDWL[428] LDWL[427]
+ LDWL[426] LDWL[425] LDWL[424] LDWL[423] LDWL[422] LDWL[421] LDWL[420] LDWL[419] LDWL[418] LDWL[417] LDWL[416]
+ LDWL[415] LDWL[414] LDWL[413] LDWL[412] LDWL[411] LDWL[410] LDWL[409] LDWL[408] LDWL[407] LDWL[406] LDWL[405]
+ LDWL[404] LDWL[403] LDWL[402] LDWL[401] LDWL[400] LDWL[399] LDWL[398] LDWL[397] LDWL[396] LDWL[395] LDWL[394]
+ LDWL[393] LDWL[392] LDWL[391] LDWL[390] LDWL[389] LDWL[388] LDWL[387] LDWL[386] LDWL[385] LDWL[384] LDWL[383]
+ LDWL[382] LDWL[381] LDWL[380] LDWL[379] LDWL[378] LDWL[377] LDWL[376] LDWL[375] LDWL[374] LDWL[373] LDWL[372]
+ LDWL[371] LDWL[370] LDWL[369] LDWL[368] LDWL[367] LDWL[366] LDWL[365] LDWL[364] LDWL[363] LDWL[362] LDWL[361]
+ LDWL[360] LDWL[359] LDWL[358] LDWL[357] LDWL[356] LDWL[355] LDWL[354] LDWL[353] LDWL[352] LDWL[351] LDWL[350]
+ LDWL[349] LDWL[348] LDWL[347] LDWL[346] LDWL[345] LDWL[344] LDWL[343] LDWL[342] LDWL[341] LDWL[340] LDWL[339]
+ LDWL[338] LDWL[337] LDWL[336] LDWL[335] LDWL[334] LDWL[333] LDWL[332] LDWL[331] LDWL[330] LDWL[329] LDWL[328]
+ LDWL[327] LDWL[326] LDWL[325] LDWL[324] LDWL[323] LDWL[322] LDWL[321] LDWL[320] LDWL[319] LDWL[318] LDWL[317]
+ LDWL[316] LDWL[315] LDWL[314] LDWL[313] LDWL[312] LDWL[311] LDWL[310] LDWL[309] LDWL[308] LDWL[307] LDWL[306]
+ LDWL[305] LDWL[304] LDWL[303] LDWL[302] LDWL[301] LDWL[300] LDWL[299] LDWL[298] LDWL[297] LDWL[296] LDWL[295]
+ LDWL[294] LDWL[293] LDWL[292] LDWL[291] LDWL[290] LDWL[289] LDWL[288] LDWL[287] LDWL[286] LDWL[285] LDWL[284]
+ LDWL[283] LDWL[282] LDWL[281] LDWL[280] LDWL[279] LDWL[278] LDWL[277] LDWL[276] LDWL[275] LDWL[274] LDWL[273]
+ LDWL[272] LDWL[271] LDWL[270] LDWL[269] LDWL[268] LDWL[267] LDWL[266] LDWL[265] LDWL[264] LDWL[263] LDWL[262]
+ LDWL[261] LDWL[260] LDWL[259] LDWL[258] LDWL[257] LDWL[256] LDWL[255] LDWL[254] LDWL[253] LDWL[252] LDWL[251]
+ LDWL[250] LDWL[249] LDWL[248] LDWL[247] LDWL[246] LDWL[245] LDWL[244] LDWL[243] LDWL[242] LDWL[241] LDWL[240]
+ LDWL[239] LDWL[238] LDWL[237] LDWL[236] LDWL[235] LDWL[234] LDWL[233] LDWL[232] LDWL[231] LDWL[230] LDWL[229]
+ LDWL[228] LDWL[227] LDWL[226] LDWL[225] LDWL[224] LDWL[223] LDWL[222] LDWL[221] LDWL[220] LDWL[219] LDWL[218]
+ LDWL[217] LDWL[216] LDWL[215] LDWL[214] LDWL[213] LDWL[212] LDWL[211] LDWL[210] LDWL[209] LDWL[208] LDWL[207]
+ LDWL[206] LDWL[205] LDWL[204] LDWL[203] LDWL[202] LDWL[201] LDWL[200] LDWL[199] LDWL[198] LDWL[197] LDWL[196]
+ LDWL[195] LDWL[194] LDWL[193] LDWL[192] LDWL[191] LDWL[190] LDWL[189] LDWL[188] LDWL[187] LDWL[186] LDWL[185]
+ LDWL[184] LDWL[183] LDWL[182] LDWL[181] LDWL[180] LDWL[179] LDWL[178] LDWL[177] LDWL[176] LDWL[175] LDWL[174]
+ LDWL[173] LDWL[172] LDWL[171] LDWL[170] LDWL[169] LDWL[168] LDWL[167] LDWL[166] LDWL[165] LDWL[164] LDWL[163]
+ LDWL[162] LDWL[161] LDWL[160] LDWL[159] LDWL[158] LDWL[157] LDWL[156] LDWL[155] LDWL[154] LDWL[153] LDWL[152]
+ LDWL[151] LDWL[150] LDWL[149] LDWL[148] LDWL[147] LDWL[146] LDWL[145] LDWL[144] LDWL[143] LDWL[142] LDWL[141]
+ LDWL[140] LDWL[139] LDWL[138] LDWL[137] LDWL[136] LDWL[135] LDWL[134] LDWL[133] LDWL[132] LDWL[131] LDWL[130]
+ LDWL[129] LDWL[128] LDWL[127] LDWL[126] LDWL[125] LDWL[124] LDWL[123] LDWL[122] LDWL[121] LDWL[120] LDWL[119]
+ LDWL[118] LDWL[117] LDWL[116] LDWL[115] LDWL[114] LDWL[113] LDWL[112] LDWL[111] LDWL[110] LDWL[109] LDWL[108]
+ LDWL[107] LDWL[106] LDWL[105] LDWL[104] LDWL[103] LDWL[102] LDWL[101] LDWL[100] LDWL[99] LDWL[98] LDWL[97]
+ LDWL[96] LDWL[95] LDWL[94] LDWL[93] LDWL[92] LDWL[91] LDWL[90] LDWL[89] LDWL[88] LDWL[87] LDWL[86] LDWL[85]
+ LDWL[84] LDWL[83] LDWL[82] LDWL[81] LDWL[80] LDWL[79] LDWL[78] LDWL[77] LDWL[76] LDWL[75] LDWL[74] LDWL[73]
+ LDWL[72] LDWL[71] LDWL[70] LDWL[69] LDWL[68] LDWL[67] LDWL[66] LDWL[65] LDWL[64] LDWL[63] LDWL[62] LDWL[61]
+ LDWL[60] LDWL[59] LDWL[58] LDWL[57] LDWL[56] LDWL[55] LDWL[54] LDWL[53] LDWL[52] LDWL[51] LDWL[50] LDWL[49]
+ LDWL[48] LDWL[47] LDWL[46] LDWL[45] LDWL[44] LDWL[43] LDWL[42] LDWL[41] LDWL[40] LDWL[39] LDWL[38] LDWL[37]
+ LDWL[36] LDWL[35] LDWL[34] LDWL[33] LDWL[32] LDWL[31] LDWL[30] LDWL[29] LDWL[28] LDWL[27] LDWL[26] LDWL[25]
+ LDWL[24] LDWL[23] LDWL[22] LDWL[21] LDWL[20] LDWL[19] LDWL[18] LDWL[17] LDWL[16] LDWL[15] LDWL[14] LDWL[13]
+ LDWL[12] LDWL[11] LDWL[10] LDWL[9] LDWL[8] LDWL[7] LDWL[6] LDWL[5] LDWL[4] LDWL[3] LDWL[2] LDWL[1] LDWL[0]
+ LDBL[255] LDBL[254] LDBL[253] LDBL[252] LDBL[251] LDBL[250] LDBL[249] LDBL[248] LDBL[247] LDBL[246] LDBL[245]
+ LDBL[244] LDBL[243] LDBL[242] LDBL[241] LDBL[240] LDBL[239] LDBL[238] LDBL[237] LDBL[236] LDBL[235] LDBL[234]
+ LDBL[233] LDBL[232] LDBL[231] LDBL[230] LDBL[229] LDBL[228] LDBL[227] LDBL[226] LDBL[225] LDBL[224] LDBL[223]
+ LDBL[222] LDBL[221] LDBL[220] LDBL[219] LDBL[218] LDBL[217] LDBL[216] LDBL[215] LDBL[214] LDBL[213] LDBL[212]
+ LDBL[211] LDBL[210] LDBL[209] LDBL[208] LDBL[207] LDBL[206] LDBL[205] LDBL[204] LDBL[203] LDBL[202] LDBL[201]
+ LDBL[200] LDBL[199] LDBL[198] LDBL[197] LDBL[196] LDBL[195] LDBL[194] LDBL[193] LDBL[192] LDBL[191] LDBL[190]
+ LDBL[189] LDBL[188] LDBL[187] LDBL[186] LDBL[185] LDBL[184] LDBL[183] LDBL[182] LDBL[181] LDBL[180] LDBL[179]
+ LDBL[178] LDBL[177] LDBL[176] LDBL[175] LDBL[174] LDBL[173] LDBL[172] LDBL[171] LDBL[170] LDBL[169] LDBL[168]
+ LDBL[167] LDBL[166] LDBL[165] LDBL[164] LDBL[163] LDBL[162] LDBL[161] LDBL[160] LDBL[159] LDBL[158] LDBL[157]
+ LDBL[156] LDBL[155] LDBL[154] LDBL[153] LDBL[152] LDBL[151] LDBL[150] LDBL[149] LDBL[148] LDBL[147] LDBL[146]
+ LDBL[145] LDBL[144] LDBL[143] LDBL[142] LDBL[141] LDBL[140] LDBL[139] LDBL[138] LDBL[137] LDBL[136] LDBL[135]
+ LDBL[134] LDBL[133] LDBL[132] LDBL[131] LDBL[130] LDBL[129] LDBL[128] LDBL[127] LDBL[126] LDBL[125] LDBL[124]
+ LDBL[123] LDBL[122] LDBL[121] LDBL[120] LDBL[119] LDBL[118] LDBL[117] LDBL[116] LDBL[115] LDBL[114] LDBL[113]
+ LDBL[112] LDBL[111] LDBL[110] LDBL[109] LDBL[108] LDBL[107] LDBL[106] LDBL[105] LDBL[104] LDBL[103] LDBL[102]
+ LDBL[101] LDBL[100] LDBL[99] LDBL[98] LDBL[97] LDBL[96] LDBL[95] LDBL[94] LDBL[93] LDBL[92] LDBL[91] LDBL[90]
+ LDBL[89] LDBL[88] LDBL[87] LDBL[86] LDBL[85] LDBL[84] LDBL[83] LDBL[82] LDBL[81] LDBL[80] LDBL[79] LDBL[78]
+ LDBL[77] LDBL[76] LDBL[75] LDBL[74] LDBL[73] LDBL[72] LDBL[71] LDBL[70] LDBL[69] LDBL[68] LDBL[67] LDBL[66]
+ LDBL[65] LDBL[64] LDBL[63] LDBL[62] LDBL[61] LDBL[60] LDBL[59] LDBL[58] LDBL[57] LDBL[56] LDBL[55] LDBL[54]
+ LDBL[53] LDBL[52] LDBL[51] LDBL[50] LDBL[49] LDBL[48] LDBL[47] LDBL[46] LDBL[45] LDBL[44] LDBL[43] LDBL[42]
+ LDBL[41] LDBL[40] LDBL[39] LDBL[38] LDBL[37] LDBL[36] LDBL[35] LDBL[34] LDBL[33] LDBL[32] LDBL[31] LDBL[30]
+ LDBL[29] LDBL[28] LDBL[27] LDBL[26] LDBL[25] LDBL[24] LDBL[23] LDBL[22] LDBL[21] LDBL[20] LDBL[19] LDBL[18]
+ LDBL[17] LDBL[16] LDBL[15] LDBL[14] LDBL[13] LDBL[12] LDBL[11] LDBL[10] LDBL[9] LDBL[8] LDBL[7] LDBL[6]
+ LDBL[5] LDBL[4] LDBL[3] LDBL[2] LDBL[1] LDBL[0] vss
*.ipin
*+ LDWL[511],LDWL[510],LDWL[509],LDWL[508],LDWL[507],LDWL[506],LDWL[505],LDWL[504],LDWL[503],LDWL[502],LDWL[501],LDWL[500],LDWL[499],LDWL[498],LDWL[497],LDWL[496],LDWL[495],LDWL[494],LDWL[493],LDWL[492],LDWL[491],LDWL[490],LDWL[489],LDWL[488],LDWL[487],LDWL[486],LDWL[485],LDWL[484],LDWL[483],LDWL[482],LDWL[481],LDWL[480],LDWL[479],LDWL[478],LDWL[477],LDWL[476],LDWL[475],LDWL[474],LDWL[473],LDWL[472],LDWL[471],LDWL[470],LDWL[469],LDWL[468],LDWL[467],LDWL[466],LDWL[465],LDWL[464],LDWL[463],LDWL[462],LDWL[461],LDWL[460],LDWL[459],LDWL[458],LDWL[457],LDWL[456],LDWL[455],LDWL[454],LDWL[453],LDWL[452],LDWL[451],LDWL[450],LDWL[449],LDWL[448],LDWL[447],LDWL[446],LDWL[445],LDWL[444],LDWL[443],LDWL[442],LDWL[441],LDWL[440],LDWL[439],LDWL[438],LDWL[437],LDWL[436],LDWL[435],LDWL[434],LDWL[433],LDWL[432],LDWL[431],LDWL[430],LDWL[429],LDWL[428],LDWL[427],LDWL[426],LDWL[425],LDWL[424],LDWL[423],LDWL[422],LDWL[421],LDWL[420],LDWL[419],LDWL[418],LDWL[417],LDWL[416],LDWL[415],LDWL[414],LDWL[413],LDWL[412],LDWL[411],LDWL[410],LDWL[409],LDWL[408],LDWL[407],LDWL[406],LDWL[405],LDWL[404],LDWL[403],LDWL[402],LDWL[401],LDWL[400],LDWL[399],LDWL[398],LDWL[397],LDWL[396],LDWL[395],LDWL[394],LDWL[393],LDWL[392],LDWL[391],LDWL[390],LDWL[389],LDWL[388],LDWL[387],LDWL[386],LDWL[385],LDWL[384],LDWL[383],LDWL[382],LDWL[381],LDWL[380],LDWL[379],LDWL[378],LDWL[377],LDWL[376],LDWL[375],LDWL[374],LDWL[373],LDWL[372],LDWL[371],LDWL[370],LDWL[369],LDWL[368],LDWL[367],LDWL[366],LDWL[365],LDWL[364],LDWL[363],LDWL[362],LDWL[361],LDWL[360],LDWL[359],LDWL[358],LDWL[357],LDWL[356],LDWL[355],LDWL[354],LDWL[353],LDWL[352],LDWL[351],LDWL[350],LDWL[349],LDWL[348],LDWL[347],LDWL[346],LDWL[345],LDWL[344],LDWL[343],LDWL[342],LDWL[341],LDWL[340],LDWL[339],LDWL[338],LDWL[337],LDWL[336],LDWL[335],LDWL[334],LDWL[333],LDWL[332],LDWL[331],LDWL[330],LDWL[329],LDWL[328],LDWL[327],LDWL[326],LDWL[325],LDWL[324],LDWL[323],LDWL[322],LDWL[321],LDWL[320],LDWL[319],LDWL[318],LDWL[317],LDWL[316],LDWL[315],LDWL[314],LDWL[313],LDWL[312],LDWL[311],LDWL[310],LDWL[309],LDWL[308],LDWL[307],LDWL[306],LDWL[305],LDWL[304],LDWL[303],LDWL[302],LDWL[301],LDWL[300],LDWL[299],LDWL[298],LDWL[297],LDWL[296],LDWL[295],LDWL[294],LDWL[293],LDWL[292],LDWL[291],LDWL[290],LDWL[289],LDWL[288],LDWL[287],LDWL[286],LDWL[285],LDWL[284],LDWL[283],LDWL[282],LDWL[281],LDWL[280],LDWL[279],LDWL[278],LDWL[277],LDWL[276],LDWL[275],LDWL[274],LDWL[273],LDWL[272],LDWL[271],LDWL[270],LDWL[269],LDWL[268],LDWL[267],LDWL[266],LDWL[265],LDWL[264],LDWL[263],LDWL[262],LDWL[261],LDWL[260],LDWL[259],LDWL[258],LDWL[257],LDWL[256],LDWL[255],LDWL[254],LDWL[253],LDWL[252],LDWL[251],LDWL[250],LDWL[249],LDWL[248],LDWL[247],LDWL[246],LDWL[245],LDWL[244],LDWL[243],LDWL[242],LDWL[241],LDWL[240],LDWL[239],LDWL[238],LDWL[237],LDWL[236],LDWL[235],LDWL[234],LDWL[233],LDWL[232],LDWL[231],LDWL[230],LDWL[229],LDWL[228],LDWL[227],LDWL[226],LDWL[225],LDWL[224],LDWL[223],LDWL[222],LDWL[221],LDWL[220],LDWL[219],LDWL[218],LDWL[217],LDWL[216],LDWL[215],LDWL[214],LDWL[213],LDWL[212],LDWL[211],LDWL[210],LDWL[209],LDWL[208],LDWL[207],LDWL[206],LDWL[205],LDWL[204],LDWL[203],LDWL[202],LDWL[201],LDWL[200],LDWL[199],LDWL[198],LDWL[197],LDWL[196],LDWL[195],LDWL[194],LDWL[193],LDWL[192],LDWL[191],LDWL[190],LDWL[189],LDWL[188],LDWL[187],LDWL[186],LDWL[185],LDWL[184],LDWL[183],LDWL[182],LDWL[181],LDWL[180],LDWL[179],LDWL[178],LDWL[177],LDWL[176],LDWL[175],LDWL[174],LDWL[173],LDWL[172],LDWL[171],LDWL[170],LDWL[169],LDWL[168],LDWL[167],LDWL[166],LDWL[165],LDWL[164],LDWL[163],LDWL[162],LDWL[161],LDWL[160],LDWL[159],LDWL[158],LDWL[157],LDWL[156],LDWL[155],LDWL[154],LDWL[153],LDWL[152],LDWL[151],LDWL[150],LDWL[149],LDWL[148],LDWL[147],LDWL[146],LDWL[145],LDWL[144],LDWL[143],LDWL[142],LDWL[141],LDWL[140],LDWL[139],LDWL[138],LDWL[137],LDWL[136],LDWL[135],LDWL[134],LDWL[133],LDWL[132],LDWL[131],LDWL[130],LDWL[129],LDWL[128],LDWL[127],LDWL[126],LDWL[125],LDWL[124],LDWL[123],LDWL[122],LDWL[121],LDWL[120],LDWL[119],LDWL[118],LDWL[117],LDWL[116],LDWL[115],LDWL[114],LDWL[113],LDWL[112],LDWL[111],LDWL[110],LDWL[109],LDWL[108],LDWL[107],LDWL[106],LDWL[105],LDWL[104],LDWL[103],LDWL[102],LDWL[101],LDWL[100],LDWL[99],LDWL[98],LDWL[97],LDWL[96],LDWL[95],LDWL[94],LDWL[93],LDWL[92],LDWL[91],LDWL[90],LDWL[89],LDWL[88],LDWL[87],LDWL[86],LDWL[85],LDWL[84],LDWL[83],LDWL[82],LDWL[81],LDWL[80],LDWL[79],LDWL[78],LDWL[77],LDWL[76],LDWL[75],LDWL[74],LDWL[73],LDWL[72],LDWL[71],LDWL[70],LDWL[69],LDWL[68],LDWL[67],LDWL[66],LDWL[65],LDWL[64],LDWL[63],LDWL[62],LDWL[61],LDWL[60],LDWL[59],LDWL[58],LDWL[57],LDWL[56],LDWL[55],LDWL[54],LDWL[53],LDWL[52],LDWL[51],LDWL[50],LDWL[49],LDWL[48],LDWL[47],LDWL[46],LDWL[45],LDWL[44],LDWL[43],LDWL[42],LDWL[41],LDWL[40],LDWL[39],LDWL[38],LDWL[37],LDWL[36],LDWL[35],LDWL[34],LDWL[33],LDWL[32],LDWL[31],LDWL[30],LDWL[29],LDWL[28],LDWL[27],LDWL[26],LDWL[25],LDWL[24],LDWL[23],LDWL[22],LDWL[21],LDWL[20],LDWL[19],LDWL[18],LDWL[17],LDWL[16],LDWL[15],LDWL[14],LDWL[13],LDWL[12],LDWL[11],LDWL[10],LDWL[9],LDWL[8],LDWL[7],LDWL[6],LDWL[5],LDWL[4],LDWL[3],LDWL[2],LDWL[1],LDWL[0]
*.iopin
*+ LDBL[255],LDBL[254],LDBL[253],LDBL[252],LDBL[251],LDBL[250],LDBL[249],LDBL[248],LDBL[247],LDBL[246],LDBL[245],LDBL[244],LDBL[243],LDBL[242],LDBL[241],LDBL[240],LDBL[239],LDBL[238],LDBL[237],LDBL[236],LDBL[235],LDBL[234],LDBL[233],LDBL[232],LDBL[231],LDBL[230],LDBL[229],LDBL[228],LDBL[227],LDBL[226],LDBL[225],LDBL[224],LDBL[223],LDBL[222],LDBL[221],LDBL[220],LDBL[219],LDBL[218],LDBL[217],LDBL[216],LDBL[215],LDBL[214],LDBL[213],LDBL[212],LDBL[211],LDBL[210],LDBL[209],LDBL[208],LDBL[207],LDBL[206],LDBL[205],LDBL[204],LDBL[203],LDBL[202],LDBL[201],LDBL[200],LDBL[199],LDBL[198],LDBL[197],LDBL[196],LDBL[195],LDBL[194],LDBL[193],LDBL[192],LDBL[191],LDBL[190],LDBL[189],LDBL[188],LDBL[187],LDBL[186],LDBL[185],LDBL[184],LDBL[183],LDBL[182],LDBL[181],LDBL[180],LDBL[179],LDBL[178],LDBL[177],LDBL[176],LDBL[175],LDBL[174],LDBL[173],LDBL[172],LDBL[171],LDBL[170],LDBL[169],LDBL[168],LDBL[167],LDBL[166],LDBL[165],LDBL[164],LDBL[163],LDBL[162],LDBL[161],LDBL[160],LDBL[159],LDBL[158],LDBL[157],LDBL[156],LDBL[155],LDBL[154],LDBL[153],LDBL[152],LDBL[151],LDBL[150],LDBL[149],LDBL[148],LDBL[147],LDBL[146],LDBL[145],LDBL[144],LDBL[143],LDBL[142],LDBL[141],LDBL[140],LDBL[139],LDBL[138],LDBL[137],LDBL[136],LDBL[135],LDBL[134],LDBL[133],LDBL[132],LDBL[131],LDBL[130],LDBL[129],LDBL[128],LDBL[127],LDBL[126],LDBL[125],LDBL[124],LDBL[123],LDBL[122],LDBL[121],LDBL[120],LDBL[119],LDBL[118],LDBL[117],LDBL[116],LDBL[115],LDBL[114],LDBL[113],LDBL[112],LDBL[111],LDBL[110],LDBL[109],LDBL[108],LDBL[107],LDBL[106],LDBL[105],LDBL[104],LDBL[103],LDBL[102],LDBL[101],LDBL[100],LDBL[99],LDBL[98],LDBL[97],LDBL[96],LDBL[95],LDBL[94],LDBL[93],LDBL[92],LDBL[91],LDBL[90],LDBL[89],LDBL[88],LDBL[87],LDBL[86],LDBL[85],LDBL[84],LDBL[83],LDBL[82],LDBL[81],LDBL[80],LDBL[79],LDBL[78],LDBL[77],LDBL[76],LDBL[75],LDBL[74],LDBL[73],LDBL[72],LDBL[71],LDBL[70],LDBL[69],LDBL[68],LDBL[67],LDBL[66],LDBL[65],LDBL[64],LDBL[63],LDBL[62],LDBL[61],LDBL[60],LDBL[59],LDBL[58],LDBL[57],LDBL[56],LDBL[55],LDBL[54],LDBL[53],LDBL[52],LDBL[51],LDBL[50],LDBL[49],LDBL[48],LDBL[47],LDBL[46],LDBL[45],LDBL[44],LDBL[43],LDBL[42],LDBL[41],LDBL[40],LDBL[39],LDBL[38],LDBL[37],LDBL[36],LDBL[35],LDBL[34],LDBL[33],LDBL[32],LDBL[31],LDBL[30],LDBL[29],LDBL[28],LDBL[27],LDBL[26],LDBL[25],LDBL[24],LDBL[23],LDBL[22],LDBL[21],LDBL[20],LDBL[19],LDBL[18],LDBL[17],LDBL[16],LDBL[15],LDBL[14],LDBL[13],LDBL[12],LDBL[11],LDBL[10],LDBL[9],LDBL[8],LDBL[7],LDBL[6],LDBL[5],LDBL[4],LDBL[3],LDBL[2],LDBL[1],LDBL[0]
*.ipin vss
c1[255] LDBL[255] 0 180f m=1
c1[254] LDBL[254] 0 180f m=1
c1[253] LDBL[253] 0 180f m=1
c1[252] LDBL[252] 0 180f m=1
c1[251] LDBL[251] 0 180f m=1
c1[250] LDBL[250] 0 180f m=1
c1[249] LDBL[249] 0 180f m=1
c1[248] LDBL[248] 0 180f m=1
c1[247] LDBL[247] 0 180f m=1
c1[246] LDBL[246] 0 180f m=1
c1[245] LDBL[245] 0 180f m=1
c1[244] LDBL[244] 0 180f m=1
c1[243] LDBL[243] 0 180f m=1
c1[242] LDBL[242] 0 180f m=1
c1[241] LDBL[241] 0 180f m=1
c1[240] LDBL[240] 0 180f m=1
c1[239] LDBL[239] 0 180f m=1
c1[238] LDBL[238] 0 180f m=1
c1[237] LDBL[237] 0 180f m=1
c1[236] LDBL[236] 0 180f m=1
c1[235] LDBL[235] 0 180f m=1
c1[234] LDBL[234] 0 180f m=1
c1[233] LDBL[233] 0 180f m=1
c1[232] LDBL[232] 0 180f m=1
c1[231] LDBL[231] 0 180f m=1
c1[230] LDBL[230] 0 180f m=1
c1[229] LDBL[229] 0 180f m=1
c1[228] LDBL[228] 0 180f m=1
c1[227] LDBL[227] 0 180f m=1
c1[226] LDBL[226] 0 180f m=1
c1[225] LDBL[225] 0 180f m=1
c1[224] LDBL[224] 0 180f m=1
c1[223] LDBL[223] 0 180f m=1
c1[222] LDBL[222] 0 180f m=1
c1[221] LDBL[221] 0 180f m=1
c1[220] LDBL[220] 0 180f m=1
c1[219] LDBL[219] 0 180f m=1
c1[218] LDBL[218] 0 180f m=1
c1[217] LDBL[217] 0 180f m=1
c1[216] LDBL[216] 0 180f m=1
c1[215] LDBL[215] 0 180f m=1
c1[214] LDBL[214] 0 180f m=1
c1[213] LDBL[213] 0 180f m=1
c1[212] LDBL[212] 0 180f m=1
c1[211] LDBL[211] 0 180f m=1
c1[210] LDBL[210] 0 180f m=1
c1[209] LDBL[209] 0 180f m=1
c1[208] LDBL[208] 0 180f m=1
c1[207] LDBL[207] 0 180f m=1
c1[206] LDBL[206] 0 180f m=1
c1[205] LDBL[205] 0 180f m=1
c1[204] LDBL[204] 0 180f m=1
c1[203] LDBL[203] 0 180f m=1
c1[202] LDBL[202] 0 180f m=1
c1[201] LDBL[201] 0 180f m=1
c1[200] LDBL[200] 0 180f m=1
c1[199] LDBL[199] 0 180f m=1
c1[198] LDBL[198] 0 180f m=1
c1[197] LDBL[197] 0 180f m=1
c1[196] LDBL[196] 0 180f m=1
c1[195] LDBL[195] 0 180f m=1
c1[194] LDBL[194] 0 180f m=1
c1[193] LDBL[193] 0 180f m=1
c1[192] LDBL[192] 0 180f m=1
c1[191] LDBL[191] 0 180f m=1
c1[190] LDBL[190] 0 180f m=1
c1[189] LDBL[189] 0 180f m=1
c1[188] LDBL[188] 0 180f m=1
c1[187] LDBL[187] 0 180f m=1
c1[186] LDBL[186] 0 180f m=1
c1[185] LDBL[185] 0 180f m=1
c1[184] LDBL[184] 0 180f m=1
c1[183] LDBL[183] 0 180f m=1
c1[182] LDBL[182] 0 180f m=1
c1[181] LDBL[181] 0 180f m=1
c1[180] LDBL[180] 0 180f m=1
c1[179] LDBL[179] 0 180f m=1
c1[178] LDBL[178] 0 180f m=1
c1[177] LDBL[177] 0 180f m=1
c1[176] LDBL[176] 0 180f m=1
c1[175] LDBL[175] 0 180f m=1
c1[174] LDBL[174] 0 180f m=1
c1[173] LDBL[173] 0 180f m=1
c1[172] LDBL[172] 0 180f m=1
c1[171] LDBL[171] 0 180f m=1
c1[170] LDBL[170] 0 180f m=1
c1[169] LDBL[169] 0 180f m=1
c1[168] LDBL[168] 0 180f m=1
c1[167] LDBL[167] 0 180f m=1
c1[166] LDBL[166] 0 180f m=1
c1[165] LDBL[165] 0 180f m=1
c1[164] LDBL[164] 0 180f m=1
c1[163] LDBL[163] 0 180f m=1
c1[162] LDBL[162] 0 180f m=1
c1[161] LDBL[161] 0 180f m=1
c1[160] LDBL[160] 0 180f m=1
c1[159] LDBL[159] 0 180f m=1
c1[158] LDBL[158] 0 180f m=1
c1[157] LDBL[157] 0 180f m=1
c1[156] LDBL[156] 0 180f m=1
c1[155] LDBL[155] 0 180f m=1
c1[154] LDBL[154] 0 180f m=1
c1[153] LDBL[153] 0 180f m=1
c1[152] LDBL[152] 0 180f m=1
c1[151] LDBL[151] 0 180f m=1
c1[150] LDBL[150] 0 180f m=1
c1[149] LDBL[149] 0 180f m=1
c1[148] LDBL[148] 0 180f m=1
c1[147] LDBL[147] 0 180f m=1
c1[146] LDBL[146] 0 180f m=1
c1[145] LDBL[145] 0 180f m=1
c1[144] LDBL[144] 0 180f m=1
c1[143] LDBL[143] 0 180f m=1
c1[142] LDBL[142] 0 180f m=1
c1[141] LDBL[141] 0 180f m=1
c1[140] LDBL[140] 0 180f m=1
c1[139] LDBL[139] 0 180f m=1
c1[138] LDBL[138] 0 180f m=1
c1[137] LDBL[137] 0 180f m=1
c1[136] LDBL[136] 0 180f m=1
c1[135] LDBL[135] 0 180f m=1
c1[134] LDBL[134] 0 180f m=1
c1[133] LDBL[133] 0 180f m=1
c1[132] LDBL[132] 0 180f m=1
c1[131] LDBL[131] 0 180f m=1
c1[130] LDBL[130] 0 180f m=1
c1[129] LDBL[129] 0 180f m=1
c1[128] LDBL[128] 0 180f m=1
c1[127] LDBL[127] 0 180f m=1
c1[126] LDBL[126] 0 180f m=1
c1[125] LDBL[125] 0 180f m=1
c1[124] LDBL[124] 0 180f m=1
c1[123] LDBL[123] 0 180f m=1
c1[122] LDBL[122] 0 180f m=1
c1[121] LDBL[121] 0 180f m=1
c1[120] LDBL[120] 0 180f m=1
c1[119] LDBL[119] 0 180f m=1
c1[118] LDBL[118] 0 180f m=1
c1[117] LDBL[117] 0 180f m=1
c1[116] LDBL[116] 0 180f m=1
c1[115] LDBL[115] 0 180f m=1
c1[114] LDBL[114] 0 180f m=1
c1[113] LDBL[113] 0 180f m=1
c1[112] LDBL[112] 0 180f m=1
c1[111] LDBL[111] 0 180f m=1
c1[110] LDBL[110] 0 180f m=1
c1[109] LDBL[109] 0 180f m=1
c1[108] LDBL[108] 0 180f m=1
c1[107] LDBL[107] 0 180f m=1
c1[106] LDBL[106] 0 180f m=1
c1[105] LDBL[105] 0 180f m=1
c1[104] LDBL[104] 0 180f m=1
c1[103] LDBL[103] 0 180f m=1
c1[102] LDBL[102] 0 180f m=1
c1[101] LDBL[101] 0 180f m=1
c1[100] LDBL[100] 0 180f m=1
c1[99] LDBL[99] 0 180f m=1
c1[98] LDBL[98] 0 180f m=1
c1[97] LDBL[97] 0 180f m=1
c1[96] LDBL[96] 0 180f m=1
c1[95] LDBL[95] 0 180f m=1
c1[94] LDBL[94] 0 180f m=1
c1[93] LDBL[93] 0 180f m=1
c1[92] LDBL[92] 0 180f m=1
c1[91] LDBL[91] 0 180f m=1
c1[90] LDBL[90] 0 180f m=1
c1[89] LDBL[89] 0 180f m=1
c1[88] LDBL[88] 0 180f m=1
c1[87] LDBL[87] 0 180f m=1
c1[86] LDBL[86] 0 180f m=1
c1[85] LDBL[85] 0 180f m=1
c1[84] LDBL[84] 0 180f m=1
c1[83] LDBL[83] 0 180f m=1
c1[82] LDBL[82] 0 180f m=1
c1[81] LDBL[81] 0 180f m=1
c1[80] LDBL[80] 0 180f m=1
c1[79] LDBL[79] 0 180f m=1
c1[78] LDBL[78] 0 180f m=1
c1[77] LDBL[77] 0 180f m=1
c1[76] LDBL[76] 0 180f m=1
c1[75] LDBL[75] 0 180f m=1
c1[74] LDBL[74] 0 180f m=1
c1[73] LDBL[73] 0 180f m=1
c1[72] LDBL[72] 0 180f m=1
c1[71] LDBL[71] 0 180f m=1
c1[70] LDBL[70] 0 180f m=1
c1[69] LDBL[69] 0 180f m=1
c1[68] LDBL[68] 0 180f m=1
c1[67] LDBL[67] 0 180f m=1
c1[66] LDBL[66] 0 180f m=1
c1[65] LDBL[65] 0 180f m=1
c1[64] LDBL[64] 0 180f m=1
c1[63] LDBL[63] 0 180f m=1
c1[62] LDBL[62] 0 180f m=1
c1[61] LDBL[61] 0 180f m=1
c1[60] LDBL[60] 0 180f m=1
c1[59] LDBL[59] 0 180f m=1
c1[58] LDBL[58] 0 180f m=1
c1[57] LDBL[57] 0 180f m=1
c1[56] LDBL[56] 0 180f m=1
c1[55] LDBL[55] 0 180f m=1
c1[54] LDBL[54] 0 180f m=1
c1[53] LDBL[53] 0 180f m=1
c1[52] LDBL[52] 0 180f m=1
c1[51] LDBL[51] 0 180f m=1
c1[50] LDBL[50] 0 180f m=1
c1[49] LDBL[49] 0 180f m=1
c1[48] LDBL[48] 0 180f m=1
c1[47] LDBL[47] 0 180f m=1
c1[46] LDBL[46] 0 180f m=1
c1[45] LDBL[45] 0 180f m=1
c1[44] LDBL[44] 0 180f m=1
c1[43] LDBL[43] 0 180f m=1
c1[42] LDBL[42] 0 180f m=1
c1[41] LDBL[41] 0 180f m=1
c1[40] LDBL[40] 0 180f m=1
c1[39] LDBL[39] 0 180f m=1
c1[38] LDBL[38] 0 180f m=1
c1[37] LDBL[37] 0 180f m=1
c1[36] LDBL[36] 0 180f m=1
c1[35] LDBL[35] 0 180f m=1
c1[34] LDBL[34] 0 180f m=1
c1[33] LDBL[33] 0 180f m=1
c1[32] LDBL[32] 0 180f m=1
c1[31] LDBL[31] 0 180f m=1
c1[30] LDBL[30] 0 180f m=1
c1[29] LDBL[29] 0 180f m=1
c1[28] LDBL[28] 0 180f m=1
c1[27] LDBL[27] 0 180f m=1
c1[26] LDBL[26] 0 180f m=1
c1[25] LDBL[25] 0 180f m=1
c1[24] LDBL[24] 0 180f m=1
c1[23] LDBL[23] 0 180f m=1
c1[22] LDBL[22] 0 180f m=1
c1[21] LDBL[21] 0 180f m=1
c1[20] LDBL[20] 0 180f m=1
c1[19] LDBL[19] 0 180f m=1
c1[18] LDBL[18] 0 180f m=1
c1[17] LDBL[17] 0 180f m=1
c1[16] LDBL[16] 0 180f m=1
c1[15] LDBL[15] 0 180f m=1
c1[14] LDBL[14] 0 180f m=1
c1[13] LDBL[13] 0 180f m=1
c1[12] LDBL[12] 0 180f m=1
c1[11] LDBL[11] 0 180f m=1
c1[10] LDBL[10] 0 180f m=1
c1[9] LDBL[9] 0 180f m=1
c1[8] LDBL[8] 0 180f m=1
c1[7] LDBL[7] 0 180f m=1
c1[6] LDBL[6] 0 180f m=1
c1[5] LDBL[5] 0 180f m=1
c1[4] LDBL[4] 0 180f m=1
c1[3] LDBL[3] 0 180f m=1
c1[2] LDBL[2] 0 180f m=1
c1[1] LDBL[1] 0 180f m=1
c1[0] LDBL[0] 0 180f m=1
**** begin user architecture code
*   pattern=1a87   word=0   wl=0 address=0000
m0 LDBL[0] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m1 LDBL[16] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m2 LDBL[32] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m3 float1 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m4 float2 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m5 float3 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m6 float4 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m7 LDBL[112] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m8 float5 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m9 LDBL[144] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m10 float6 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m11 LDBL[176] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m12 LDBL[192] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m13 float7 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m14 float8 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m15 float9 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
*   pattern=0298   word=1   wl=0 address=0001
m16 float10 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m17 float11 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m18 float12 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m19 LDBL[49] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m20 LDBL[65] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m21 float13 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m22 float14 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m23 LDBL[113] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m24 float15 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m25 LDBL[145] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m26 float16 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m27 float17 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m28 float18 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m29 float19 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m30 float20 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m31 float21 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
*   pattern=aa6a   word=2   wl=0 address=0002
m32 float22 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m33 LDBL[18] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m34 float23 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m35 LDBL[50] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m36 float24 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m37 LDBL[82] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m38 LDBL[98] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m39 float25 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m40 float26 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m41 LDBL[146] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m42 float27 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m43 LDBL[178] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m44 float28 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m45 LDBL[210] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m46 float29 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m47 LDBL[242] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f719   word=3   wl=0 address=0003
m48 LDBL[3] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m49 float30 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m50 float31 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m51 LDBL[51] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m52 LDBL[67] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m53 float32 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m54 float33 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m55 float34 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m56 LDBL[131] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m57 LDBL[147] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m58 LDBL[163] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m59 float35 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m60 LDBL[195] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m61 LDBL[211] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m62 LDBL[227] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m63 LDBL[243] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=eb3e   word=4   wl=0 address=0004
m64 float36 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m65 LDBL[20] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m66 LDBL[36] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m67 LDBL[52] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m68 LDBL[68] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m69 LDBL[84] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m70 float37 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m71 float38 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m72 LDBL[132] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m73 LDBL[148] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m74 float39 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m75 LDBL[180] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m76 float40 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m77 LDBL[212] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m78 LDBL[228] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m79 LDBL[244] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4bd0   word=5   wl=0 address=0005
m80 float41 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m81 float42 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m82 float43 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m83 float44 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m84 LDBL[69] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m85 float45 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m86 LDBL[101] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m87 LDBL[117] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m88 LDBL[133] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m89 LDBL[149] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m90 float46 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m91 LDBL[181] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m92 float47 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m93 float48 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m94 LDBL[229] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m95 float49 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
*   pattern=1039   word=6   wl=0 address=0006
m96 LDBL[6] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m97 float50 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m98 float51 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m99 LDBL[54] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m100 LDBL[70] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m101 LDBL[86] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m102 float52 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m103 float53 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m104 float54 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m105 float55 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m106 float56 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m107 float57 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m108 LDBL[198] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m109 float58 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m110 float59 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m111 float60 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
*   pattern=86aa   word=7   wl=0 address=0007
m112 float61 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m113 LDBL[23] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m114 float62 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m115 LDBL[55] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m116 float63 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m117 LDBL[87] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m118 float64 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m119 LDBL[119] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m120 float65 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m121 LDBL[151] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m122 LDBL[167] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m123 float66 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m124 float67 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m125 float68 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m126 float69 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m127 LDBL[247] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b708   word=8   wl=0 address=0008
m128 float70 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m129 float71 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m130 float72 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m131 LDBL[56] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m132 float73 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m133 float74 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m134 float75 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m135 float76 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m136 LDBL[136] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m137 LDBL[152] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m138 LDBL[168] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m139 float77 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m140 LDBL[200] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m141 LDBL[216] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m142 float78 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m143 LDBL[248] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a07e   word=9   wl=0 address=0009
m144 float79 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m145 LDBL[25] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m146 LDBL[41] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m147 LDBL[57] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m148 LDBL[73] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m149 LDBL[89] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m150 LDBL[105] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m151 float80 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m152 float81 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m153 float82 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m154 float83 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m155 float84 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m156 float85 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m157 LDBL[217] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m158 float86 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m159 LDBL[249] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=13e8   word=10   wl=0 address=000a
m160 float87 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m161 float88 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m162 float89 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m163 LDBL[58] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m164 float90 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m165 LDBL[90] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m166 LDBL[106] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m167 LDBL[122] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m168 LDBL[138] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m169 LDBL[154] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m170 float91 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m171 float92 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m172 LDBL[202] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m173 float93 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m174 float94 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m175 float95 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
*   pattern=387e   word=11   wl=0 address=000b
m176 float96 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m177 LDBL[27] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m178 LDBL[43] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m179 LDBL[59] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m180 LDBL[75] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m181 LDBL[91] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m182 LDBL[107] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m183 float97 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m184 float98 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m185 float99 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m186 float100 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m187 LDBL[187] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m188 LDBL[203] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m189 LDBL[219] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m190 float101 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m191 float102 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2172   word=12   wl=0 address=000c
m192 float103 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m193 LDBL[28] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m194 float104 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m195 float105 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m196 LDBL[76] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m197 LDBL[92] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m198 LDBL[108] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m199 float106 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m200 LDBL[140] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m201 float107 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m202 float108 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m203 float109 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m204 float110 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m205 LDBL[220] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m206 float111 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m207 float112 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1553   word=13   wl=0 address=000d
m208 LDBL[13] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m209 LDBL[29] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m210 float113 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m211 float114 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m212 LDBL[77] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m213 float115 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m214 LDBL[109] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m215 float116 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m216 LDBL[141] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m217 float117 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m218 LDBL[173] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m219 float118 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m220 LDBL[205] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m221 float119 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m222 float120 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m223 float121 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=90cf   word=14   wl=0 address=000e
m224 LDBL[14] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m225 LDBL[30] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m226 LDBL[46] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m227 LDBL[62] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m228 float122 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m229 float123 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m230 LDBL[110] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m231 LDBL[126] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m232 float124 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m233 float125 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m234 float126 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m235 float127 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m236 LDBL[206] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m237 float128 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m238 float129 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m239 LDBL[254] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9c87   word=15   wl=0 address=000f
m240 LDBL[15] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m241 LDBL[31] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m242 LDBL[47] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m243 float130 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m244 float131 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m245 float132 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m246 float133 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m247 LDBL[127] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m248 float134 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m249 float135 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m250 LDBL[175] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m251 LDBL[191] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m252 LDBL[207] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m253 float136 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m254 float137 LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m255 LDBL[255] LDWL[0] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=508f   word=0   wl=1 address=0010
m256 LDBL[0] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m257 LDBL[16] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m258 LDBL[32] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m259 LDBL[48] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m260 float138 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m261 float139 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m262 float140 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m263 LDBL[112] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m264 float141 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m265 float142 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m266 float143 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m267 float144 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m268 LDBL[192] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m269 float145 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m270 LDBL[224] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m271 float146 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9bb4   word=1   wl=1 address=0011
m272 float147 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m273 float148 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m274 LDBL[33] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m275 float149 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m276 LDBL[65] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m277 LDBL[81] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m278 float150 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m279 LDBL[113] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m280 LDBL[129] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m281 LDBL[145] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m282 float151 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m283 LDBL[177] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m284 LDBL[193] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m285 float152 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m286 float153 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m287 LDBL[241] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3abb   word=2   wl=1 address=0012
m288 LDBL[2] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m289 LDBL[18] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m290 float154 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m291 LDBL[50] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m292 LDBL[66] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m293 LDBL[82] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m294 float155 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m295 LDBL[114] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m296 float156 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m297 LDBL[146] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m298 float157 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m299 LDBL[178] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m300 LDBL[194] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m301 LDBL[210] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m302 float158 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m303 float159 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c209   word=3   wl=1 address=0013
m304 LDBL[3] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m305 float160 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m306 float161 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m307 LDBL[51] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m308 float162 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m309 float163 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m310 float164 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m311 float165 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m312 float166 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m313 LDBL[147] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m314 float167 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m315 float168 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m316 float169 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m317 float170 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m318 LDBL[227] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m319 LDBL[243] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a6e9   word=4   wl=1 address=0014
m320 LDBL[4] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m321 float171 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m322 float172 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m323 LDBL[52] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m324 float173 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m325 LDBL[84] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m326 LDBL[100] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m327 LDBL[116] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m328 float174 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m329 LDBL[148] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m330 LDBL[164] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m331 float175 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m332 float176 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m333 LDBL[212] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m334 float177 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m335 LDBL[244] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a4a3   word=5   wl=1 address=0015
m336 LDBL[5] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m337 LDBL[21] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m338 float178 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m339 float179 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m340 float180 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m341 LDBL[85] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m342 float181 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m343 LDBL[117] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m344 float182 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m345 float183 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m346 LDBL[165] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m347 float184 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m348 float185 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m349 LDBL[213] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m350 float186 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m351 LDBL[245] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ac53   word=6   wl=1 address=0016
m352 LDBL[6] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m353 LDBL[22] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m354 float187 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m355 float188 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m356 LDBL[70] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m357 float189 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m358 LDBL[102] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m359 float190 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m360 float191 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m361 float192 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m362 LDBL[166] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m363 LDBL[182] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m364 float193 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m365 LDBL[214] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m366 float194 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m367 LDBL[246] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b070   word=7   wl=1 address=0017
m368 float195 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m369 float196 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m370 float197 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m371 float198 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m372 LDBL[71] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m373 LDBL[87] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m374 LDBL[103] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m375 float199 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m376 float200 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m377 float201 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m378 float202 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m379 float203 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m380 LDBL[199] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m381 LDBL[215] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m382 float204 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m383 LDBL[247] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=42fd   word=8   wl=1 address=0018
m384 LDBL[8] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m385 float205 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m386 LDBL[40] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m387 LDBL[56] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m388 LDBL[72] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m389 LDBL[88] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m390 LDBL[104] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m391 LDBL[120] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m392 float206 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m393 LDBL[152] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m394 float207 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m395 float208 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m396 float209 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m397 float210 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m398 LDBL[232] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m399 float211 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=74dd   word=9   wl=1 address=0019
m400 LDBL[9] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m401 float212 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m402 LDBL[41] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m403 LDBL[57] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m404 LDBL[73] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m405 float213 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m406 LDBL[105] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m407 LDBL[121] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m408 float214 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m409 float215 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m410 LDBL[169] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m411 float216 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m412 LDBL[201] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m413 LDBL[217] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m414 LDBL[233] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m415 float217 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6bab   word=10   wl=1 address=001a
m416 LDBL[10] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m417 LDBL[26] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m418 float218 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m419 LDBL[58] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m420 float219 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m421 LDBL[90] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m422 float220 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m423 LDBL[122] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m424 LDBL[138] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m425 LDBL[154] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m426 float221 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m427 LDBL[186] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m428 float222 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m429 LDBL[218] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m430 LDBL[234] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m431 float223 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a39a   word=11   wl=1 address=001b
m432 float224 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m433 LDBL[27] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m434 float225 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m435 LDBL[59] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m436 LDBL[75] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m437 float226 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m438 float227 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m439 LDBL[123] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m440 LDBL[139] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m441 LDBL[155] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m442 float228 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m443 float229 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m444 float230 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m445 LDBL[219] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m446 float231 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m447 LDBL[251] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2110   word=12   wl=1 address=001c
m448 float232 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m449 float233 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m450 float234 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m451 float235 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m452 LDBL[76] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m453 float236 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m454 float237 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m455 float238 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m456 LDBL[140] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m457 float239 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m458 float240 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m459 float241 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m460 float242 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m461 LDBL[220] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m462 float243 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m463 float244 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ce81   word=13   wl=1 address=001d
m464 LDBL[13] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m465 float245 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m466 float246 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m467 float247 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m468 float248 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m469 float249 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m470 float250 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m471 LDBL[125] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m472 float251 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m473 LDBL[157] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m474 LDBL[173] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m475 LDBL[189] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m476 float252 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m477 float253 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m478 LDBL[237] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m479 LDBL[253] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a021   word=14   wl=1 address=001e
m480 LDBL[14] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m481 float254 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m482 float255 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m483 float256 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m484 float257 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m485 LDBL[94] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m486 float258 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m487 float259 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m488 float260 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m489 float261 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m490 float262 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m491 float263 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m492 float264 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m493 LDBL[222] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m494 float265 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m495 LDBL[254] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ce52   word=15   wl=1 address=001f
m496 float266 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m497 LDBL[31] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m498 float267 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m499 float268 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m500 LDBL[79] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m501 float269 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m502 LDBL[111] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m503 float270 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m504 float271 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m505 LDBL[159] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m506 LDBL[175] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m507 LDBL[191] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m508 float272 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m509 float273 LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m510 LDBL[239] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m511 LDBL[255] LDWL[1] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=016e   word=0   wl=2 address=0020
m512 float274 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m513 LDBL[16] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m514 LDBL[32] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m515 LDBL[48] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m516 float275 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m517 LDBL[80] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m518 LDBL[96] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m519 float276 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m520 LDBL[128] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m521 float277 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m522 float278 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m523 float279 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m524 float280 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m525 float281 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m526 float282 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m527 float283 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=57f6   word=1   wl=2 address=0021
m528 float284 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m529 LDBL[17] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m530 LDBL[33] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m531 float285 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m532 LDBL[65] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m533 LDBL[81] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m534 LDBL[97] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m535 LDBL[113] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m536 LDBL[129] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m537 LDBL[145] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m538 LDBL[161] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m539 float286 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m540 LDBL[193] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m541 float287 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m542 LDBL[225] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m543 float288 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b835   word=2   wl=2 address=0022
m544 LDBL[2] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m545 float289 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m546 LDBL[34] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m547 float290 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m548 LDBL[66] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m549 LDBL[82] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m550 float291 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m551 float292 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m552 float293 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m553 float294 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m554 float295 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m555 LDBL[178] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m556 LDBL[194] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m557 LDBL[210] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m558 float296 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m559 LDBL[242] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=406a   word=3   wl=2 address=0023
m560 float297 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m561 LDBL[19] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m562 float298 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m563 LDBL[51] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m564 float299 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m565 LDBL[83] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m566 LDBL[99] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m567 float300 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m568 float301 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m569 float302 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m570 float303 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m571 float304 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m572 float305 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m573 float306 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m574 LDBL[227] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m575 float307 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6877   word=4   wl=2 address=0024
m576 LDBL[4] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m577 LDBL[20] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m578 LDBL[36] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m579 float308 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m580 LDBL[68] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m581 LDBL[84] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m582 LDBL[100] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m583 float309 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m584 float310 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m585 float311 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m586 float312 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m587 LDBL[180] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m588 float313 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m589 LDBL[212] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m590 LDBL[228] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m591 float314 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ace7   word=5   wl=2 address=0025
m592 LDBL[5] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m593 LDBL[21] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m594 LDBL[37] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m595 float315 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m596 float316 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m597 LDBL[85] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m598 LDBL[101] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m599 LDBL[117] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m600 float317 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m601 float318 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m602 LDBL[165] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m603 LDBL[181] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m604 float319 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m605 LDBL[213] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m606 float320 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m607 LDBL[245] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1e49   word=6   wl=2 address=0026
m608 LDBL[6] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m609 float321 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m610 float322 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m611 LDBL[54] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m612 float323 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m613 float324 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m614 LDBL[102] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m615 float325 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m616 float326 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m617 LDBL[150] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m618 LDBL[166] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m619 LDBL[182] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m620 LDBL[198] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m621 float327 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m622 float328 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m623 float329 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6c31   word=7   wl=2 address=0027
m624 LDBL[7] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m625 float330 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m626 float331 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m627 float332 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m628 LDBL[71] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m629 LDBL[87] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m630 float333 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m631 float334 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m632 float335 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m633 float336 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m634 LDBL[167] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m635 LDBL[183] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m636 float337 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m637 LDBL[215] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m638 LDBL[231] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m639 float338 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d027   word=8   wl=2 address=0028
m640 LDBL[8] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m641 LDBL[24] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m642 LDBL[40] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m643 float339 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m644 float340 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m645 LDBL[88] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m646 float341 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m647 float342 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m648 float343 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m649 float344 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m650 float345 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m651 float346 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m652 LDBL[200] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m653 float347 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m654 LDBL[232] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m655 LDBL[248] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b89b   word=9   wl=2 address=0029
m656 LDBL[9] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m657 LDBL[25] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m658 float348 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m659 LDBL[57] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m660 LDBL[73] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m661 float349 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m662 float350 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m663 LDBL[121] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m664 float351 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m665 float352 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m666 float353 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m667 LDBL[185] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m668 LDBL[201] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m669 LDBL[217] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m670 float354 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m671 LDBL[249] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fceb   word=10   wl=2 address=002a
m672 LDBL[10] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m673 LDBL[26] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m674 float355 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m675 LDBL[58] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m676 float356 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m677 LDBL[90] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m678 LDBL[106] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m679 LDBL[122] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m680 float357 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m681 float358 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m682 LDBL[170] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m683 LDBL[186] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m684 LDBL[202] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m685 LDBL[218] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m686 LDBL[234] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m687 LDBL[250] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9615   word=11   wl=2 address=002b
m688 LDBL[11] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m689 float359 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m690 LDBL[43] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m691 float360 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m692 LDBL[75] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m693 float361 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m694 float362 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m695 float363 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m696 float364 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m697 LDBL[155] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m698 LDBL[171] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m699 float365 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m700 LDBL[203] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m701 float366 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m702 float367 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m703 LDBL[251] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8723   word=12   wl=2 address=002c
m704 LDBL[12] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m705 LDBL[28] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m706 float368 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m707 float369 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m708 float370 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m709 LDBL[92] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m710 float371 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m711 float372 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m712 LDBL[140] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m713 LDBL[156] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m714 LDBL[172] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m715 float373 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m716 float374 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m717 float375 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m718 float376 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m719 LDBL[252] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=05ad   word=13   wl=2 address=002d
m720 LDBL[13] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m721 float377 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m722 LDBL[45] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m723 LDBL[61] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m724 float378 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m725 LDBL[93] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m726 float379 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m727 LDBL[125] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m728 LDBL[141] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m729 float380 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m730 LDBL[173] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m731 float381 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m732 float382 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m733 float383 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m734 float384 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m735 float385 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b9d4   word=14   wl=2 address=002e
m736 float386 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m737 float387 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m738 LDBL[46] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m739 float388 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m740 LDBL[78] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m741 float389 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m742 LDBL[110] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m743 LDBL[126] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m744 LDBL[142] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m745 float390 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m746 float391 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m747 LDBL[190] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m748 LDBL[206] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m749 LDBL[222] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m750 float392 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m751 LDBL[254] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3b7e   word=15   wl=2 address=002f
m752 float393 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m753 LDBL[31] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m754 LDBL[47] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m755 LDBL[63] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m756 LDBL[79] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m757 LDBL[95] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m758 LDBL[111] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m759 float394 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m760 LDBL[143] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m761 LDBL[159] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m762 float395 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m763 LDBL[191] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m764 LDBL[207] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m765 LDBL[223] LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m766 float396 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m767 float397 LDWL[2] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d0f0   word=0   wl=3 address=0030
m768 float398 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m769 float399 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m770 float400 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m771 float401 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m772 LDBL[64] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m773 LDBL[80] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m774 LDBL[96] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m775 LDBL[112] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m776 float402 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m777 float403 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m778 float404 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m779 float405 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m780 LDBL[192] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m781 float406 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m782 LDBL[224] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m783 LDBL[240] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=88ec   word=1   wl=3 address=0031
m784 float407 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m785 float408 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m786 LDBL[33] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m787 LDBL[49] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m788 float409 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m789 LDBL[81] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m790 LDBL[97] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m791 LDBL[113] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m792 float410 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m793 float411 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m794 float412 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m795 LDBL[177] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m796 float413 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m797 float414 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m798 float415 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m799 LDBL[241] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a62c   word=2   wl=3 address=0032
m800 float416 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m801 float417 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m802 LDBL[34] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m803 LDBL[50] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m804 float418 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m805 LDBL[82] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m806 float419 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m807 float420 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m808 float421 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m809 LDBL[146] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m810 LDBL[162] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m811 float422 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m812 float423 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m813 LDBL[210] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m814 float424 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m815 LDBL[242] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=22f4   word=3   wl=3 address=0033
m816 float425 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m817 float426 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m818 LDBL[35] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m819 float427 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m820 LDBL[67] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m821 LDBL[83] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m822 LDBL[99] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m823 LDBL[115] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m824 float428 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m825 LDBL[147] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m826 float429 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m827 float430 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m828 float431 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m829 LDBL[211] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m830 float432 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m831 float433 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5ead   word=4   wl=3 address=0034
m832 LDBL[4] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m833 float434 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m834 LDBL[36] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m835 LDBL[52] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m836 float435 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m837 LDBL[84] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m838 float436 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m839 LDBL[116] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m840 float437 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m841 LDBL[148] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m842 LDBL[164] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m843 LDBL[180] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m844 LDBL[196] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m845 float438 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m846 LDBL[228] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m847 float439 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=88ae   word=5   wl=3 address=0035
m848 float440 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m849 LDBL[21] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m850 LDBL[37] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m851 LDBL[53] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m852 float441 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m853 LDBL[85] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m854 float442 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m855 LDBL[117] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m856 float443 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m857 float444 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m858 float445 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m859 LDBL[181] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m860 float446 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m861 float447 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m862 float448 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m863 LDBL[245] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8296   word=6   wl=3 address=0036
m864 float449 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m865 LDBL[22] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m866 LDBL[38] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m867 float450 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m868 LDBL[70] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m869 float451 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m870 float452 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m871 LDBL[118] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m872 float453 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m873 LDBL[150] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m874 float454 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m875 float455 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m876 float456 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m877 float457 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m878 float458 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m879 LDBL[246] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1851   word=7   wl=3 address=0037
m880 LDBL[7] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m881 float459 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m882 float460 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m883 float461 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m884 LDBL[71] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m885 float462 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m886 LDBL[103] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m887 float463 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m888 float464 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m889 float465 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m890 float466 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m891 LDBL[183] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m892 LDBL[199] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m893 float467 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m894 float468 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m895 float469 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a961   word=8   wl=3 address=0038
m896 LDBL[8] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06 m=1
m897 float470 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m898 float471 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m899 float472 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m900 float473 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m901 LDBL[88] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m902 LDBL[104] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m903 float474 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m904 LDBL[136] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m905 float475 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m906 float476 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m907 LDBL[184] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m908 float477 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m909 LDBL[216] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m910 float478 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m911 LDBL[248] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f95c   word=9   wl=3 address=0039
m912 float479 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m913 float480 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m914 LDBL[41] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m915 LDBL[57] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m916 LDBL[73] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m917 float481 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m918 LDBL[105] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m919 float482 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m920 LDBL[137] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m921 float483 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m922 float484 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m923 LDBL[185] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m924 LDBL[201] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m925 LDBL[217] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m926 LDBL[233] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m927 LDBL[249] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=595f   word=10   wl=3 address=003a
m928 LDBL[10] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m929 LDBL[26] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m930 LDBL[42] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m931 LDBL[58] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m932 LDBL[74] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m933 float485 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m934 LDBL[106] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m935 float486 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m936 LDBL[138] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m937 float487 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m938 float488 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m939 LDBL[186] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m940 LDBL[202] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m941 float489 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m942 LDBL[234] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m943 float490 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3f07   word=11   wl=3 address=003b
m944 LDBL[11] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m945 LDBL[27] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m946 LDBL[43] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m947 float491 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m948 float492 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m949 float493 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m950 float494 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m951 float495 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m952 LDBL[139] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m953 LDBL[155] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m954 LDBL[171] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m955 LDBL[187] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m956 LDBL[203] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m957 LDBL[219] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m958 float496 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m959 float497 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a056   word=12   wl=3 address=003c
m960 float498 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m961 LDBL[28] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m962 LDBL[44] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m963 float499 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m964 LDBL[76] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m965 float500 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m966 LDBL[108] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m967 float501 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m968 float502 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m969 float503 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m970 float504 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m971 float505 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m972 float506 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m973 LDBL[220] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m974 float507 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m975 LDBL[252] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9200   word=13   wl=3 address=003d
m976 float508 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m977 float509 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m978 float510 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m979 float511 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m980 float512 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m981 float513 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m982 float514 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m983 float515 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m984 float516 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m985 LDBL[157] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m986 float517 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m987 float518 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m988 LDBL[205] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m989 float519 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m990 float520 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m991 LDBL[253] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4a9f   word=14   wl=3 address=003e
m992 LDBL[14] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m993 LDBL[30] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m994 LDBL[46] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m995 LDBL[62] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m996 LDBL[78] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m997 float521 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m998 float522 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m999 LDBL[126] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1000 float523 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1001 LDBL[158] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1002 float524 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1003 LDBL[190] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1004 float525 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1005 float526 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1006 LDBL[238] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1007 float527 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=14ff   word=15   wl=3 address=003f
m1008 LDBL[15] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1009 LDBL[31] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1010 LDBL[47] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1011 LDBL[63] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1012 LDBL[79] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1013 LDBL[95] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1014 LDBL[111] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1015 LDBL[127] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1016 float528 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1017 float529 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1018 LDBL[175] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1019 float530 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1020 LDBL[207] LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1021 float531 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1022 float532 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1023 float533 LDWL[3] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1419   word=0   wl=4 address=0040
m1024 LDBL[0] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1025 float534 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1026 float535 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1027 LDBL[48] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1028 LDBL[64] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1029 float536 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1030 float537 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1031 float538 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1032 float539 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1033 float540 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1034 LDBL[160] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1035 float541 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1036 LDBL[192] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1037 float542 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1038 float543 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1039 float544 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=98b6   word=1   wl=4 address=0041
m1040 float545 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1041 LDBL[17] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1042 LDBL[33] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1043 float546 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1044 LDBL[65] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1045 LDBL[81] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1046 float547 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1047 LDBL[113] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1048 float548 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1049 float549 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1050 float550 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1051 LDBL[177] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1052 LDBL[193] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1053 float551 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1054 float552 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1055 LDBL[241] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9c4b   word=2   wl=4 address=0042
m1056 LDBL[2] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1057 LDBL[18] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1058 float553 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1059 LDBL[50] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1060 float554 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1061 float555 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1062 LDBL[98] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1063 float556 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1064 float557 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1065 float558 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1066 LDBL[162] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1067 LDBL[178] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1068 LDBL[194] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1069 float559 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1070 float560 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1071 LDBL[242] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8fc2   word=3   wl=4 address=0043
m1072 float561 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1073 LDBL[19] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1074 float562 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1075 float563 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1076 float564 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1077 float565 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1078 LDBL[99] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1079 LDBL[115] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1080 LDBL[131] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1081 LDBL[147] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1082 LDBL[163] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1083 LDBL[179] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1084 float566 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1085 float567 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1086 float568 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1087 LDBL[243] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=bb4f   word=4   wl=4 address=0044
m1088 LDBL[4] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1089 LDBL[20] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1090 LDBL[36] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1091 LDBL[52] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1092 float569 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1093 float570 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1094 LDBL[100] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1095 float571 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1096 LDBL[132] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1097 LDBL[148] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1098 float572 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1099 LDBL[180] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1100 LDBL[196] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1101 LDBL[212] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1102 float573 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1103 LDBL[244] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c0cd   word=5   wl=4 address=0045
m1104 LDBL[5] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1105 float574 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1106 LDBL[37] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1107 LDBL[53] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1108 float575 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1109 float576 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1110 LDBL[101] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1111 LDBL[117] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1112 float577 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1113 float578 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1114 float579 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1115 float580 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1116 float581 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1117 float582 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1118 LDBL[229] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1119 LDBL[245] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=06aa   word=6   wl=4 address=0046
m1120 float583 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1121 LDBL[22] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1122 float584 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1123 LDBL[54] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1124 float585 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1125 LDBL[86] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1126 float586 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1127 LDBL[118] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1128 float587 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1129 LDBL[150] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1130 LDBL[166] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1131 float588 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1132 float589 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1133 float590 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1134 float591 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1135 float592 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3dd8   word=7   wl=4 address=0047
m1136 float593 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1137 float594 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1138 float595 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1139 LDBL[55] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1140 LDBL[71] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1141 float596 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1142 LDBL[103] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1143 LDBL[119] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1144 LDBL[135] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1145 float597 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1146 LDBL[167] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1147 LDBL[183] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1148 LDBL[199] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1149 LDBL[215] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1150 float598 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1151 float599 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=52da   word=8   wl=4 address=0048
m1152 float600 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1153 LDBL[24] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1154 float601 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1155 LDBL[56] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1156 LDBL[72] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1157 float602 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1158 LDBL[104] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1159 LDBL[120] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1160 float603 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1161 LDBL[152] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1162 float604 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1163 float605 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1164 LDBL[200] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1165 float606 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1166 LDBL[232] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1167 float607 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=be0b   word=9   wl=4 address=0049
m1168 LDBL[9] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1169 LDBL[25] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1170 float608 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1171 LDBL[57] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1172 float609 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1173 float610 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1174 float611 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1175 float612 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1176 float613 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1177 LDBL[153] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1178 LDBL[169] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1179 LDBL[185] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1180 LDBL[201] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1181 LDBL[217] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1182 float614 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1183 LDBL[249] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f912   word=10   wl=4 address=004a
m1184 float615 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1185 LDBL[26] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1186 float616 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1187 float617 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1188 LDBL[74] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1189 float618 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1190 float619 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1191 float620 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1192 LDBL[138] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1193 float621 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1194 float622 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1195 LDBL[186] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1196 LDBL[202] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1197 LDBL[218] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1198 LDBL[234] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1199 LDBL[250] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4edc   word=11   wl=4 address=004b
m1200 float623 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1201 float624 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1202 LDBL[43] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1203 LDBL[59] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1204 LDBL[75] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1205 float625 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1206 LDBL[107] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1207 LDBL[123] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1208 float626 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1209 LDBL[155] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1210 LDBL[171] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1211 LDBL[187] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1212 float627 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1213 float628 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1214 LDBL[235] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1215 float629 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9d40   word=12   wl=4 address=004c
m1216 float630 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1217 float631 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1218 float632 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1219 float633 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1220 float634 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1221 float635 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1222 LDBL[108] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1223 float636 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1224 LDBL[140] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1225 float637 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1226 LDBL[172] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1227 LDBL[188] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1228 LDBL[204] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1229 float638 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1230 float639 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1231 LDBL[252] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2ef0   word=13   wl=4 address=004d
m1232 float640 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1233 float641 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1234 float642 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1235 float643 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1236 LDBL[77] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1237 LDBL[93] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1238 LDBL[109] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1239 LDBL[125] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1240 float644 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1241 LDBL[157] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1242 LDBL[173] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1243 LDBL[189] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1244 float645 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1245 LDBL[221] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1246 float646 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1247 float647 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c914   word=14   wl=4 address=004e
m1248 float648 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1249 float649 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1250 LDBL[46] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1251 float650 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1252 LDBL[78] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1253 float651 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1254 float652 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1255 float653 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1256 LDBL[142] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1257 float654 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1258 float655 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1259 LDBL[190] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1260 float656 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1261 float657 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1262 LDBL[238] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1263 LDBL[254] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fe34   word=15   wl=4 address=004f
m1264 float658 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1265 float659 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1266 LDBL[47] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1267 float660 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1268 LDBL[79] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1269 LDBL[95] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1270 float661 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1271 float662 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1272 float663 LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1273 LDBL[159] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1274 LDBL[175] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1275 LDBL[191] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1276 LDBL[207] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1277 LDBL[223] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1278 LDBL[239] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1279 LDBL[255] LDWL[4] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=837d   word=0   wl=5 address=0050
m1280 LDBL[0] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1281 float664 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1282 LDBL[32] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1283 LDBL[48] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1284 LDBL[64] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1285 LDBL[80] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1286 LDBL[96] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1287 float665 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1288 LDBL[128] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1289 LDBL[144] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1290 float666 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1291 float667 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1292 float668 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1293 float669 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1294 float670 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1295 LDBL[240] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e2c4   word=1   wl=5 address=0051
m1296 float671 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1297 float672 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1298 LDBL[33] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1299 float673 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1300 float674 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1301 float675 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1302 LDBL[97] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1303 LDBL[113] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1304 float676 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1305 LDBL[145] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1306 float677 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1307 float678 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1308 float679 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1309 LDBL[209] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1310 LDBL[225] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1311 LDBL[241] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c133   word=2   wl=5 address=0052
m1312 LDBL[2] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1313 LDBL[18] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1314 float680 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1315 float681 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1316 LDBL[66] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1317 LDBL[82] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1318 float682 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1319 float683 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1320 LDBL[130] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1321 float684 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1322 float685 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1323 float686 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1324 float687 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1325 float688 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1326 LDBL[226] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1327 LDBL[242] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=53d8   word=3   wl=5 address=0053
m1328 float689 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1329 float690 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1330 float691 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1331 LDBL[51] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1332 LDBL[67] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1333 float692 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1334 LDBL[99] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1335 LDBL[115] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1336 LDBL[131] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1337 LDBL[147] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1338 float693 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1339 float694 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1340 LDBL[195] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1341 float695 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1342 LDBL[227] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1343 float696 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8b92   word=4   wl=5 address=0054
m1344 float697 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1345 LDBL[20] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1346 float698 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1347 float699 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1348 LDBL[68] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1349 float700 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1350 float701 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1351 LDBL[116] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1352 LDBL[132] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1353 LDBL[148] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1354 float702 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1355 LDBL[180] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1356 float703 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1357 float704 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1358 float705 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1359 LDBL[244] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=54ec   word=5   wl=5 address=0055
m1360 float706 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1361 float707 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1362 LDBL[37] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1363 LDBL[53] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1364 float708 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1365 LDBL[85] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1366 LDBL[101] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1367 LDBL[117] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1368 float709 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1369 float710 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1370 LDBL[165] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1371 float711 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1372 LDBL[197] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1373 float712 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1374 LDBL[229] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1375 float713 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9aa7   word=6   wl=5 address=0056
m1376 LDBL[6] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1377 LDBL[22] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1378 LDBL[38] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1379 float714 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1380 float715 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1381 LDBL[86] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1382 float716 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1383 LDBL[118] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1384 float717 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1385 LDBL[150] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1386 float718 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1387 LDBL[182] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1388 LDBL[198] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1389 float719 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1390 float720 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1391 LDBL[246] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=add8   word=7   wl=5 address=0057
m1392 float721 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1393 float722 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1394 float723 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1395 LDBL[55] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1396 LDBL[71] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1397 float724 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1398 LDBL[103] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1399 LDBL[119] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1400 LDBL[135] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1401 float725 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1402 LDBL[167] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1403 LDBL[183] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1404 float726 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1405 LDBL[215] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1406 float727 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1407 LDBL[247] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=34b4   word=8   wl=5 address=0058
m1408 float728 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1409 float729 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1410 LDBL[40] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1411 float730 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1412 LDBL[72] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1413 LDBL[88] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1414 float731 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1415 LDBL[120] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1416 float732 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1417 float733 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1418 LDBL[168] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1419 float734 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1420 LDBL[200] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1421 LDBL[216] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1422 float735 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1423 float736 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6e5c   word=9   wl=5 address=0059
m1424 float737 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1425 float738 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1426 LDBL[41] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1427 LDBL[57] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1428 LDBL[73] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1429 float739 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1430 LDBL[105] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1431 float740 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1432 float741 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1433 LDBL[153] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1434 LDBL[169] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1435 LDBL[185] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1436 float742 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1437 LDBL[217] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1438 LDBL[233] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1439 float743 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c464   word=10   wl=5 address=005a
m1440 float744 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1441 float745 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1442 LDBL[42] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1443 float746 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1444 float747 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1445 LDBL[90] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1446 LDBL[106] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1447 float748 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1448 float749 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1449 float750 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1450 LDBL[170] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1451 float751 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1452 float752 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1453 float753 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1454 LDBL[234] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1455 LDBL[250] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=35a5   word=11   wl=5 address=005b
m1456 LDBL[11] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1457 float754 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1458 LDBL[43] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1459 float755 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1460 float756 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1461 LDBL[91] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1462 float757 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1463 LDBL[123] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1464 LDBL[139] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1465 float758 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1466 LDBL[171] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1467 float759 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1468 LDBL[203] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1469 LDBL[219] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1470 float760 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1471 float761 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4a4b   word=12   wl=5 address=005c
m1472 LDBL[12] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1473 LDBL[28] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1474 float762 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1475 LDBL[60] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1476 float763 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1477 float764 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1478 LDBL[108] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1479 float765 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1480 float766 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1481 LDBL[156] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1482 float767 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1483 LDBL[188] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1484 float768 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1485 float769 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1486 LDBL[236] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1487 float770 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3458   word=13   wl=5 address=005d
m1488 float771 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1489 float772 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1490 float773 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1491 LDBL[61] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1492 LDBL[77] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1493 float774 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1494 LDBL[109] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1495 float775 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1496 float776 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1497 float777 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1498 LDBL[173] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1499 float778 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1500 LDBL[205] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1501 LDBL[221] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1502 float779 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1503 float780 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e801   word=14   wl=5 address=005e
m1504 LDBL[14] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1505 float781 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1506 float782 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1507 float783 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1508 float784 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1509 float785 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1510 float786 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1511 float787 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1512 float788 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1513 float789 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1514 float790 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1515 LDBL[190] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1516 float791 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1517 LDBL[222] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1518 LDBL[238] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1519 LDBL[254] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3451   word=15   wl=5 address=005f
m1520 LDBL[15] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1521 float792 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1522 float793 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1523 float794 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1524 LDBL[79] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1525 float795 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1526 LDBL[111] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1527 float796 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1528 float797 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1529 float798 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1530 LDBL[175] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1531 float799 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1532 LDBL[207] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1533 LDBL[223] LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1534 float800 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1535 float801 LDWL[5] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=196e   word=0   wl=6 address=0060
m1536 float802 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1537 LDBL[16] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1538 LDBL[32] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1539 LDBL[48] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1540 float803 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1541 LDBL[80] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1542 LDBL[96] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1543 float804 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1544 LDBL[128] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1545 float805 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1546 float806 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1547 LDBL[176] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1548 LDBL[192] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1549 float807 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1550 float808 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1551 float809 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=78b0   word=1   wl=6 address=0061
m1552 float810 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1553 float811 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1554 float812 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1555 float813 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1556 LDBL[65] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1557 LDBL[81] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1558 float814 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1559 LDBL[113] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1560 float815 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1561 float816 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1562 float817 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1563 LDBL[177] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1564 LDBL[193] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1565 LDBL[209] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1566 LDBL[225] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1567 float818 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=df82   word=2   wl=6 address=0062
m1568 float819 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1569 LDBL[18] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1570 float820 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1571 float821 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1572 float822 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1573 float823 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1574 float824 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1575 LDBL[114] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1576 LDBL[130] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1577 LDBL[146] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1578 LDBL[162] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1579 LDBL[178] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1580 LDBL[194] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1581 float825 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1582 LDBL[226] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1583 LDBL[242] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=139c   word=3   wl=6 address=0063
m1584 float826 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1585 float827 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1586 LDBL[35] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1587 LDBL[51] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1588 LDBL[67] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1589 float828 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1590 float829 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1591 LDBL[115] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1592 LDBL[131] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1593 LDBL[147] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1594 float830 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1595 float831 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1596 LDBL[195] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1597 float832 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1598 float833 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1599 float834 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2d17   word=4   wl=6 address=0064
m1600 LDBL[4] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1601 LDBL[20] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1602 LDBL[36] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1603 float835 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1604 LDBL[68] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1605 float836 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1606 float837 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1607 float838 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1608 LDBL[132] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1609 float839 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1610 LDBL[164] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1611 LDBL[180] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1612 float840 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1613 LDBL[212] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1614 float841 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1615 float842 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2b93   word=5   wl=6 address=0065
m1616 LDBL[5] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1617 LDBL[21] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1618 float843 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1619 float844 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1620 LDBL[69] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1621 float845 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1622 float846 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1623 LDBL[117] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1624 LDBL[133] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1625 LDBL[149] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1626 float847 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1627 LDBL[181] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1628 float848 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1629 LDBL[213] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1630 float849 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1631 float850 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=265b   word=6   wl=6 address=0066
m1632 LDBL[6] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1633 LDBL[22] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1634 float851 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1635 LDBL[54] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1636 LDBL[70] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1637 float852 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1638 LDBL[102] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1639 float853 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1640 float854 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1641 LDBL[150] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1642 LDBL[166] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1643 float855 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1644 float856 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1645 LDBL[214] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1646 float857 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1647 float858 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e7af   word=7   wl=6 address=0067
m1648 LDBL[7] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1649 LDBL[23] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1650 LDBL[39] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1651 LDBL[55] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1652 float859 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1653 LDBL[87] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1654 float860 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1655 LDBL[119] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1656 LDBL[135] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1657 LDBL[151] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1658 LDBL[167] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1659 float861 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1660 float862 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1661 LDBL[215] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1662 LDBL[231] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1663 LDBL[247] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7851   word=8   wl=6 address=0068
m1664 LDBL[8] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1665 float863 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1666 float864 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1667 float865 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1668 LDBL[72] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1669 float866 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1670 LDBL[104] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1671 float867 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1672 float868 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1673 float869 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1674 float870 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1675 LDBL[184] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1676 LDBL[200] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1677 LDBL[216] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1678 LDBL[232] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1679 float871 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=259f   word=9   wl=6 address=0069
m1680 LDBL[9] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1681 LDBL[25] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1682 LDBL[41] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1683 LDBL[57] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1684 LDBL[73] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1685 float872 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1686 float873 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1687 LDBL[121] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1688 LDBL[137] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1689 float874 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1690 LDBL[169] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1691 float875 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1692 float876 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1693 LDBL[217] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1694 float877 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1695 float878 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=94f6   word=10   wl=6 address=006a
m1696 float879 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1697 LDBL[26] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1698 LDBL[42] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1699 float880 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1700 LDBL[74] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1701 LDBL[90] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1702 LDBL[106] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1703 LDBL[122] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1704 float881 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1705 float882 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1706 LDBL[170] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1707 float883 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1708 LDBL[202] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1709 float884 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1710 float885 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1711 LDBL[250] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=764b   word=11   wl=6 address=006b
m1712 LDBL[11] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1713 LDBL[27] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1714 float886 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1715 LDBL[59] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1716 float887 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1717 float888 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1718 LDBL[107] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1719 float889 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1720 float890 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1721 LDBL[155] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1722 LDBL[171] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1723 float891 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1724 LDBL[203] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1725 LDBL[219] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1726 LDBL[235] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1727 float892 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4481   word=12   wl=6 address=006c
m1728 LDBL[12] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1729 float893 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1730 float894 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1731 float895 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1732 float896 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1733 float897 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1734 float898 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1735 LDBL[124] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1736 float899 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1737 float900 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1738 LDBL[172] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1739 float901 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1740 float902 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1741 float903 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1742 LDBL[236] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1743 float904 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3bdd   word=13   wl=6 address=006d
m1744 LDBL[13] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1745 float905 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1746 LDBL[45] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1747 LDBL[61] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1748 LDBL[77] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1749 float906 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1750 LDBL[109] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1751 LDBL[125] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1752 LDBL[141] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1753 LDBL[157] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1754 float907 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1755 LDBL[189] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1756 LDBL[205] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1757 LDBL[221] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1758 float908 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1759 float909 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7507   word=14   wl=6 address=006e
m1760 LDBL[14] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1761 LDBL[30] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1762 LDBL[46] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1763 float910 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1764 float911 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1765 float912 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1766 float913 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1767 float914 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1768 LDBL[142] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1769 float915 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1770 LDBL[174] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1771 float916 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1772 LDBL[206] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1773 LDBL[222] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1774 LDBL[238] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1775 float917 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=396e   word=15   wl=6 address=006f
m1776 float918 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1777 LDBL[31] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1778 LDBL[47] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1779 LDBL[63] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1780 float919 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1781 LDBL[95] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1782 LDBL[111] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1783 float920 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1784 LDBL[143] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1785 float921 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1786 float922 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1787 LDBL[191] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1788 LDBL[207] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1789 LDBL[223] LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1790 float923 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1791 float924 LDWL[6] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=703a   word=0   wl=7 address=0070
m1792 float925 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1793 LDBL[16] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1794 float926 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1795 LDBL[48] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1796 LDBL[64] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1797 LDBL[80] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1798 float927 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1799 float928 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1800 float929 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1801 float930 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1802 float931 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1803 float932 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1804 LDBL[192] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1805 LDBL[208] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1806 LDBL[224] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1807 float933 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f5d5   word=1   wl=7 address=0071
m1808 LDBL[1] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1809 float934 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1810 LDBL[33] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1811 float935 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1812 LDBL[65] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1813 float936 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1814 LDBL[97] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1815 LDBL[113] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1816 LDBL[129] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1817 float937 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1818 LDBL[161] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1819 float938 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1820 LDBL[193] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1821 LDBL[209] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1822 LDBL[225] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1823 LDBL[241] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1791   word=2   wl=7 address=0072
m1824 LDBL[2] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1825 float939 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1826 float940 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1827 float941 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1828 LDBL[66] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1829 float942 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1830 float943 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1831 LDBL[114] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1832 LDBL[130] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1833 LDBL[146] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1834 LDBL[162] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1835 float944 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1836 LDBL[194] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1837 float945 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1838 float946 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1839 float947 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=371c   word=3   wl=7 address=0073
m1840 float948 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1841 float949 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1842 LDBL[35] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1843 LDBL[51] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1844 LDBL[67] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1845 float950 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1846 float951 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1847 float952 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1848 LDBL[131] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1849 LDBL[147] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1850 LDBL[163] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1851 float953 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1852 LDBL[195] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1853 LDBL[211] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1854 float954 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1855 float955 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4dff   word=4   wl=7 address=0074
m1856 LDBL[4] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1857 LDBL[20] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1858 LDBL[36] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1859 LDBL[52] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1860 LDBL[68] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1861 LDBL[84] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1862 LDBL[100] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1863 LDBL[116] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1864 LDBL[132] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1865 float956 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1866 LDBL[164] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1867 LDBL[180] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1868 float957 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1869 float958 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1870 LDBL[228] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1871 float959 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3911   word=5   wl=7 address=0075
m1872 LDBL[5] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1873 float960 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1874 float961 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1875 float962 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1876 LDBL[69] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1877 float963 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1878 float964 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1879 float965 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1880 LDBL[133] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1881 float966 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1882 float967 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1883 LDBL[181] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1884 LDBL[197] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1885 LDBL[213] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1886 float968 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1887 float969 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a23a   word=6   wl=7 address=0076
m1888 float970 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1889 LDBL[22] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1890 float971 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1891 LDBL[54] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1892 LDBL[70] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1893 LDBL[86] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1894 float972 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1895 float973 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1896 float974 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1897 LDBL[150] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1898 float975 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1899 float976 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1900 float977 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1901 LDBL[214] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1902 float978 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1903 LDBL[246] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f5eb   word=7   wl=7 address=0077
m1904 LDBL[7] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1905 LDBL[23] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1906 float979 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1907 LDBL[55] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1908 float980 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1909 LDBL[87] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1910 LDBL[103] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1911 LDBL[119] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1912 LDBL[135] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1913 float981 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1914 LDBL[167] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1915 float982 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1916 LDBL[199] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1917 LDBL[215] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1918 LDBL[231] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1919 LDBL[247] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d75e   word=8   wl=7 address=0078
m1920 float983 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1921 LDBL[24] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1922 LDBL[40] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1923 LDBL[56] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1924 LDBL[72] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1925 float984 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1926 LDBL[104] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1927 float985 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1928 LDBL[136] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1929 LDBL[152] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1930 LDBL[168] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1931 float986 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1932 LDBL[200] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1933 float987 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1934 LDBL[232] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1935 LDBL[248] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2965   word=9   wl=7 address=0079
m1936 LDBL[9] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1937 float988 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1938 LDBL[41] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1939 float989 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1940 float990 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1941 LDBL[89] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1942 LDBL[105] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1943 float991 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1944 LDBL[137] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1945 float992 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1946 float993 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1947 LDBL[185] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1948 float994 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1949 LDBL[217] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1950 float995 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1951 float996 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6aaa   word=10   wl=7 address=007a
m1952 float997 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1953 LDBL[26] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1954 float998 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1955 LDBL[58] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1956 float999 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1957 LDBL[90] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1958 float1000 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1959 LDBL[122] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1960 float1001 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1961 LDBL[154] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1962 float1002 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1963 LDBL[186] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1964 float1003 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1965 LDBL[218] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1966 LDBL[234] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1967 float1004 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ec5f   word=11   wl=7 address=007b
m1968 LDBL[11] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1969 LDBL[27] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1970 LDBL[43] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1971 LDBL[59] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1972 LDBL[75] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1973 float1005 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1974 LDBL[107] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1975 float1006 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1976 float1007 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1977 float1008 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1978 LDBL[171] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1979 LDBL[187] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1980 float1009 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1981 LDBL[219] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1982 LDBL[235] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1983 LDBL[251] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a5a0   word=12   wl=7 address=007c
m1984 float1010 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1985 float1011 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1986 float1012 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1987 float1013 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1988 float1014 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1989 LDBL[92] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1990 float1015 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1991 LDBL[124] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1992 LDBL[140] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1993 float1016 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1994 LDBL[172] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1995 float1017 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1996 float1018 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1997 LDBL[220] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1998 float1019 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m1999 LDBL[252] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5ad8   word=13   wl=7 address=007d
m2000 float1020 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2001 float1021 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2002 float1022 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2003 LDBL[61] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2004 LDBL[77] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2005 float1023 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2006 LDBL[109] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2007 LDBL[125] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2008 float1024 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2009 LDBL[157] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2010 float1025 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2011 LDBL[189] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2012 LDBL[205] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2013 float1026 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2014 LDBL[237] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2015 float1027 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e317   word=14   wl=7 address=007e
m2016 LDBL[14] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2017 LDBL[30] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2018 LDBL[46] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2019 float1028 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2020 LDBL[78] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2021 float1029 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2022 float1030 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2023 float1031 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2024 LDBL[142] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2025 LDBL[158] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2026 float1032 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2027 float1033 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2028 float1034 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2029 LDBL[222] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2030 LDBL[238] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2031 LDBL[254] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3973   word=15   wl=7 address=007f
m2032 LDBL[15] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2033 LDBL[31] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2034 float1035 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2035 float1036 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2036 LDBL[79] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2037 LDBL[95] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2038 LDBL[111] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2039 float1037 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2040 LDBL[143] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2041 float1038 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2042 float1039 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2043 LDBL[191] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2044 LDBL[207] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2045 LDBL[223] LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2046 float1040 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2047 float1041 LDWL[7] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c933   word=0   wl=8 address=0080
m2048 LDBL[0] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2049 LDBL[16] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2050 float1042 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2051 float1043 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2052 LDBL[64] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2053 LDBL[80] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2054 float1044 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2055 float1045 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2056 LDBL[128] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2057 float1046 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2058 float1047 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2059 LDBL[176] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2060 float1048 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2061 float1049 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2062 LDBL[224] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2063 LDBL[240] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5164   word=1   wl=8 address=0081
m2064 float1050 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2065 float1051 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2066 LDBL[33] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2067 float1052 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2068 float1053 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2069 LDBL[81] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2070 LDBL[97] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2071 float1054 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2072 LDBL[129] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2073 float1055 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2074 float1056 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2075 float1057 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2076 LDBL[193] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2077 float1058 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2078 LDBL[225] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2079 float1059 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=115d   word=2   wl=8 address=0082
m2080 LDBL[2] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2081 float1060 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2082 LDBL[34] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2083 LDBL[50] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2084 LDBL[66] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2085 float1061 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2086 LDBL[98] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2087 float1062 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2088 LDBL[130] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2089 float1063 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2090 float1064 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2091 float1065 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2092 LDBL[194] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2093 float1066 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2094 float1067 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2095 float1068 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6a22   word=3   wl=8 address=0083
m2096 float1069 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2097 LDBL[19] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2098 float1070 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2099 float1071 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2100 float1072 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2101 LDBL[83] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2102 float1073 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2103 float1074 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2104 float1075 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2105 LDBL[147] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2106 float1076 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2107 LDBL[179] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2108 float1077 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2109 LDBL[211] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2110 LDBL[227] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2111 float1078 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8416   word=4   wl=8 address=0084
m2112 float1079 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2113 LDBL[20] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2114 LDBL[36] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2115 float1080 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2116 LDBL[68] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2117 float1081 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2118 float1082 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2119 float1083 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2120 float1084 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2121 float1085 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2122 LDBL[164] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2123 float1086 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2124 float1087 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2125 float1088 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2126 float1089 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2127 LDBL[244] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=66a4   word=5   wl=8 address=0085
m2128 float1090 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2129 float1091 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2130 LDBL[37] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2131 float1092 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2132 float1093 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2133 LDBL[85] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2134 float1094 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2135 LDBL[117] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2136 float1095 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2137 LDBL[149] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2138 LDBL[165] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2139 float1096 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2140 float1097 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2141 LDBL[213] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2142 LDBL[229] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2143 float1098 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5c63   word=6   wl=8 address=0086
m2144 LDBL[6] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2145 LDBL[22] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2146 float1099 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2147 float1100 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2148 float1101 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2149 LDBL[86] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2150 LDBL[102] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2151 float1102 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2152 float1103 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2153 float1104 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2154 LDBL[166] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2155 LDBL[182] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2156 LDBL[198] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2157 float1105 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2158 LDBL[230] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2159 float1106 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=76e0   word=7   wl=8 address=0087
m2160 float1107 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2161 float1108 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2162 float1109 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2163 float1110 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2164 float1111 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2165 LDBL[87] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2166 LDBL[103] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2167 LDBL[119] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2168 float1112 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2169 LDBL[151] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2170 LDBL[167] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2171 float1113 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2172 LDBL[199] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2173 LDBL[215] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2174 LDBL[231] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2175 float1114 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e0d5   word=8   wl=8 address=0088
m2176 LDBL[8] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2177 float1115 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2178 LDBL[40] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2179 float1116 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2180 LDBL[72] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2181 float1117 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2182 LDBL[104] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2183 LDBL[120] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2184 float1118 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2185 float1119 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2186 float1120 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2187 float1121 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2188 float1122 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2189 LDBL[216] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2190 LDBL[232] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2191 LDBL[248] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=77a5   word=9   wl=8 address=0089
m2192 LDBL[9] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2193 float1123 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2194 LDBL[41] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2195 float1124 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2196 float1125 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2197 LDBL[89] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2198 float1126 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2199 LDBL[121] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2200 LDBL[137] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2201 LDBL[153] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2202 LDBL[169] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2203 float1127 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2204 LDBL[201] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2205 LDBL[217] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2206 LDBL[233] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2207 float1128 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c4a2   word=10   wl=8 address=008a
m2208 float1129 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2209 LDBL[26] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2210 float1130 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2211 float1131 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2212 float1132 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2213 LDBL[90] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2214 float1133 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2215 LDBL[122] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2216 float1134 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2217 float1135 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2218 LDBL[170] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2219 float1136 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2220 float1137 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2221 float1138 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2222 LDBL[234] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2223 LDBL[250] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=483e   word=11   wl=8 address=008b
m2224 float1139 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2225 LDBL[27] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2226 LDBL[43] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2227 LDBL[59] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2228 LDBL[75] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2229 LDBL[91] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2230 float1140 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2231 float1141 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2232 float1142 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2233 float1143 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2234 float1144 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2235 LDBL[187] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2236 float1145 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2237 float1146 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2238 LDBL[235] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2239 float1147 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=589c   word=12   wl=8 address=008c
m2240 float1148 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2241 float1149 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2242 LDBL[44] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2243 LDBL[60] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2244 LDBL[76] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2245 float1150 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2246 float1151 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2247 LDBL[124] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2248 float1152 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2249 float1153 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2250 float1154 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2251 LDBL[188] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2252 LDBL[204] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2253 float1155 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2254 LDBL[236] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2255 float1156 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c9fc   word=13   wl=8 address=008d
m2256 float1157 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2257 float1158 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2258 LDBL[45] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2259 LDBL[61] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2260 LDBL[77] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2261 LDBL[93] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2262 LDBL[109] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2263 LDBL[125] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2264 LDBL[141] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2265 float1159 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2266 float1160 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2267 LDBL[189] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2268 float1161 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2269 float1162 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2270 LDBL[237] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2271 LDBL[253] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8542   word=14   wl=8 address=008e
m2272 float1163 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2273 LDBL[30] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2274 float1164 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2275 float1165 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2276 float1166 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2277 float1167 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2278 LDBL[110] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2279 float1168 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2280 LDBL[142] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2281 float1169 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2282 LDBL[174] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2283 float1170 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2284 float1171 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2285 float1172 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2286 float1173 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2287 LDBL[254] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a9dd   word=15   wl=8 address=008f
m2288 LDBL[15] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2289 float1174 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2290 LDBL[47] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2291 LDBL[63] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2292 LDBL[79] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2293 float1175 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2294 LDBL[111] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2295 LDBL[127] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2296 LDBL[143] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2297 float1176 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2298 float1177 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2299 LDBL[191] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2300 float1178 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2301 LDBL[223] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2302 float1179 LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2303 LDBL[255] LDWL[8] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3071   word=0   wl=9 address=0090
m2304 LDBL[0] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2305 float1180 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2306 float1181 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2307 float1182 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2308 LDBL[64] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2309 LDBL[80] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2310 LDBL[96] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2311 float1183 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2312 float1184 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2313 float1185 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2314 float1186 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2315 float1187 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2316 LDBL[192] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2317 LDBL[208] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2318 float1188 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2319 float1189 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7f08   word=1   wl=9 address=0091
m2320 float1190 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2321 float1191 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2322 float1192 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2323 LDBL[49] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2324 float1193 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2325 float1194 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2326 float1195 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2327 float1196 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2328 LDBL[129] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2329 LDBL[145] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2330 LDBL[161] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2331 LDBL[177] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2332 LDBL[193] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2333 LDBL[209] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2334 LDBL[225] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2335 float1197 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7687   word=2   wl=9 address=0092
m2336 LDBL[2] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2337 LDBL[18] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2338 LDBL[34] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2339 float1198 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2340 float1199 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2341 float1200 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2342 float1201 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2343 LDBL[114] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2344 float1202 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2345 LDBL[146] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2346 LDBL[162] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2347 float1203 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2348 LDBL[194] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2349 LDBL[210] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2350 LDBL[226] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2351 float1204 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=cbd3   word=3   wl=9 address=0093
m2352 LDBL[3] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2353 LDBL[19] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2354 float1205 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2355 float1206 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2356 LDBL[67] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2357 float1207 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2358 LDBL[99] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2359 LDBL[115] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2360 LDBL[131] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2361 LDBL[147] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2362 float1208 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2363 LDBL[179] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2364 float1209 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2365 float1210 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2366 LDBL[227] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2367 LDBL[243] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d96c   word=4   wl=9 address=0094
m2368 float1211 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2369 float1212 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2370 LDBL[36] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2371 LDBL[52] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2372 float1213 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2373 LDBL[84] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2374 LDBL[100] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2375 float1214 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2376 LDBL[132] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2377 float1215 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2378 float1216 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2379 LDBL[180] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2380 LDBL[196] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2381 float1217 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2382 LDBL[228] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2383 LDBL[244] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f6f6   word=5   wl=9 address=0095
m2384 float1218 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2385 LDBL[21] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2386 LDBL[37] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2387 float1219 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2388 LDBL[69] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2389 LDBL[85] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2390 LDBL[101] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2391 LDBL[117] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2392 float1220 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2393 LDBL[149] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2394 LDBL[165] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2395 float1221 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2396 LDBL[197] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2397 LDBL[213] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2398 LDBL[229] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2399 LDBL[245] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c9ca   word=6   wl=9 address=0096
m2400 float1222 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2401 LDBL[22] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2402 float1223 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2403 LDBL[54] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2404 float1224 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2405 float1225 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2406 LDBL[102] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2407 LDBL[118] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2408 LDBL[134] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2409 float1226 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2410 float1227 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2411 LDBL[182] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2412 float1228 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2413 float1229 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2414 LDBL[230] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2415 LDBL[246] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7f7c   word=7   wl=9 address=0097
m2416 float1230 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2417 float1231 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2418 LDBL[39] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2419 LDBL[55] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2420 LDBL[71] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2421 LDBL[87] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2422 LDBL[103] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2423 float1232 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2424 LDBL[135] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2425 LDBL[151] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2426 LDBL[167] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2427 LDBL[183] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2428 LDBL[199] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2429 LDBL[215] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2430 LDBL[231] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2431 float1233 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e714   word=8   wl=9 address=0098
m2432 float1234 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2433 float1235 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2434 LDBL[40] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2435 float1236 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2436 LDBL[72] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2437 float1237 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2438 float1238 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2439 float1239 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2440 LDBL[136] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2441 LDBL[152] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2442 LDBL[168] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2443 float1240 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2444 float1241 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2445 LDBL[216] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2446 LDBL[232] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2447 LDBL[248] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=16d2   word=9   wl=9 address=0099
m2448 float1242 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2449 LDBL[25] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2450 float1243 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2451 float1244 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2452 LDBL[73] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2453 float1245 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2454 LDBL[105] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2455 LDBL[121] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2456 float1246 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2457 LDBL[153] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2458 LDBL[169] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2459 float1247 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2460 LDBL[201] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2461 float1248 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2462 float1249 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2463 float1250 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=658d   word=10   wl=9 address=009a
m2464 LDBL[10] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2465 float1251 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2466 LDBL[42] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2467 LDBL[58] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2468 float1252 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2469 float1253 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2470 float1254 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2471 LDBL[122] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2472 LDBL[138] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2473 float1255 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2474 LDBL[170] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2475 float1256 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2476 float1257 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2477 LDBL[218] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2478 LDBL[234] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2479 float1258 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f54a   word=11   wl=9 address=009b
m2480 float1259 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2481 LDBL[27] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2482 float1260 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2483 LDBL[59] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2484 float1261 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2485 float1262 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2486 LDBL[107] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2487 float1263 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2488 LDBL[139] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2489 float1264 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2490 LDBL[171] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2491 float1265 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2492 LDBL[203] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2493 LDBL[219] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2494 LDBL[235] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2495 LDBL[251] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=acac   word=12   wl=9 address=009c
m2496 float1266 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2497 float1267 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2498 LDBL[44] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2499 LDBL[60] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2500 float1268 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2501 LDBL[92] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2502 float1269 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2503 LDBL[124] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2504 float1270 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2505 float1271 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2506 LDBL[172] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2507 LDBL[188] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2508 float1272 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2509 LDBL[220] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2510 float1273 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2511 LDBL[252] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2555   word=13   wl=9 address=009d
m2512 LDBL[13] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2513 float1274 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2514 LDBL[45] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2515 float1275 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2516 LDBL[77] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2517 float1276 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2518 LDBL[109] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2519 float1277 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2520 LDBL[141] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2521 float1278 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2522 LDBL[173] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2523 float1279 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2524 float1280 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2525 LDBL[221] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2526 float1281 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2527 float1282 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7d4f   word=14   wl=9 address=009e
m2528 LDBL[14] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2529 LDBL[30] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2530 LDBL[46] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2531 LDBL[62] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2532 float1283 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2533 float1284 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2534 LDBL[110] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2535 float1285 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2536 LDBL[142] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2537 float1286 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2538 LDBL[174] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2539 LDBL[190] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2540 LDBL[206] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2541 LDBL[222] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2542 LDBL[238] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2543 float1287 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d81b   word=15   wl=9 address=009f
m2544 LDBL[15] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2545 LDBL[31] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2546 float1288 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2547 LDBL[63] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2548 LDBL[79] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2549 float1289 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2550 float1290 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2551 float1291 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2552 float1292 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2553 float1293 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2554 float1294 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2555 LDBL[191] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2556 LDBL[207] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2557 float1295 LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2558 LDBL[239] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2559 LDBL[255] LDWL[9] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2ff1   word=0   wl=10 address=00a0
m2560 LDBL[0] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2561 float1296 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2562 float1297 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2563 float1298 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2564 LDBL[64] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2565 LDBL[80] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2566 LDBL[96] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2567 LDBL[112] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2568 LDBL[128] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2569 LDBL[144] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2570 LDBL[160] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2571 LDBL[176] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2572 float1299 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2573 LDBL[208] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2574 float1300 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2575 float1301 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=99b0   word=1   wl=10 address=00a1
m2576 float1302 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2577 float1303 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2578 float1304 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2579 float1305 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2580 LDBL[65] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2581 LDBL[81] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2582 float1306 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2583 LDBL[113] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2584 LDBL[129] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2585 float1307 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2586 float1308 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2587 LDBL[177] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2588 LDBL[193] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2589 float1309 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2590 float1310 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2591 LDBL[241] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=baae   word=2   wl=10 address=00a2
m2592 float1311 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2593 LDBL[18] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2594 LDBL[34] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2595 LDBL[50] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2596 float1312 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2597 LDBL[82] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2598 float1313 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2599 LDBL[114] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2600 float1314 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2601 LDBL[146] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2602 float1315 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2603 LDBL[178] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2604 LDBL[194] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2605 LDBL[210] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2606 float1316 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2607 LDBL[242] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0242   word=3   wl=10 address=00a3
m2608 float1317 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2609 LDBL[19] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2610 float1318 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2611 float1319 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2612 float1320 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2613 float1321 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2614 LDBL[99] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2615 float1322 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2616 float1323 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2617 LDBL[147] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2618 float1324 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2619 float1325 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2620 float1326 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2621 float1327 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2622 float1328 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2623 float1329 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=06ea   word=4   wl=10 address=00a4
m2624 float1330 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2625 LDBL[20] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2626 float1331 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2627 LDBL[52] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2628 float1332 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2629 LDBL[84] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2630 LDBL[100] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2631 LDBL[116] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2632 float1333 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2633 LDBL[148] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2634 LDBL[164] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2635 float1334 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2636 float1335 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2637 float1336 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2638 float1337 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2639 float1338 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=66f9   word=5   wl=10 address=00a5
m2640 LDBL[5] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2641 float1339 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2642 float1340 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2643 LDBL[53] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2644 LDBL[69] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2645 LDBL[85] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2646 LDBL[101] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2647 LDBL[117] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2648 float1341 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2649 LDBL[149] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2650 LDBL[165] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2651 float1342 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2652 float1343 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2653 LDBL[213] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2654 LDBL[229] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2655 float1344 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fa9a   word=6   wl=10 address=00a6
m2656 float1345 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2657 LDBL[22] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2658 float1346 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2659 LDBL[54] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2660 LDBL[70] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2661 float1347 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2662 float1348 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2663 LDBL[118] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2664 float1349 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2665 LDBL[150] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2666 float1350 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2667 LDBL[182] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2668 LDBL[198] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2669 LDBL[214] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2670 LDBL[230] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2671 LDBL[246] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=123d   word=7   wl=10 address=00a7
m2672 LDBL[7] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2673 float1351 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2674 LDBL[39] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2675 LDBL[55] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2676 LDBL[71] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2677 LDBL[87] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2678 float1352 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2679 float1353 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2680 float1354 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2681 LDBL[151] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2682 float1355 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2683 float1356 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2684 LDBL[199] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2685 float1357 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2686 float1358 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2687 float1359 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e97f   word=8   wl=10 address=00a8
m2688 LDBL[8] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2689 LDBL[24] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2690 LDBL[40] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2691 LDBL[56] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2692 LDBL[72] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2693 LDBL[88] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2694 LDBL[104] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2695 float1360 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2696 LDBL[136] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2697 float1361 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2698 float1362 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2699 LDBL[184] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2700 float1363 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2701 LDBL[216] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2702 LDBL[232] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2703 LDBL[248] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6484   word=9   wl=10 address=00a9
m2704 float1364 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2705 float1365 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2706 LDBL[41] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2707 float1366 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2708 float1367 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2709 float1368 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2710 float1369 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2711 LDBL[121] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2712 float1370 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2713 float1371 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2714 LDBL[169] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2715 float1372 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2716 float1373 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2717 LDBL[217] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2718 LDBL[233] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2719 float1374 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=19b4   word=10   wl=10 address=00aa
m2720 float1375 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2721 float1376 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2722 LDBL[42] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2723 float1377 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2724 LDBL[74] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2725 LDBL[90] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2726 float1378 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2727 LDBL[122] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2728 LDBL[138] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2729 float1379 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2730 float1380 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2731 LDBL[186] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2732 LDBL[202] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2733 float1381 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2734 float1382 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2735 float1383 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=090d   word=11   wl=10 address=00ab
m2736 LDBL[11] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2737 float1384 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2738 LDBL[43] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2739 LDBL[59] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2740 float1385 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2741 float1386 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2742 float1387 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2743 float1388 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2744 LDBL[139] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2745 float1389 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2746 float1390 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2747 LDBL[187] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2748 float1391 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2749 float1392 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2750 float1393 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2751 float1394 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8edf   word=12   wl=10 address=00ac
m2752 LDBL[12] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2753 LDBL[28] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2754 LDBL[44] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2755 LDBL[60] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2756 LDBL[76] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2757 float1395 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2758 LDBL[108] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2759 LDBL[124] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2760 float1396 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2761 LDBL[156] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2762 LDBL[172] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2763 LDBL[188] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2764 float1397 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2765 float1398 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2766 float1399 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2767 LDBL[252] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=bec6   word=13   wl=10 address=00ad
m2768 float1400 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2769 LDBL[29] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2770 LDBL[45] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2771 float1401 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2772 float1402 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2773 float1403 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2774 LDBL[109] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2775 LDBL[125] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2776 float1404 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2777 LDBL[157] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2778 LDBL[173] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2779 LDBL[189] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2780 LDBL[205] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2781 LDBL[221] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2782 float1405 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2783 LDBL[253] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7b35   word=14   wl=10 address=00ae
m2784 LDBL[14] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2785 float1406 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2786 LDBL[46] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2787 float1407 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2788 LDBL[78] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2789 LDBL[94] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2790 float1408 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2791 float1409 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2792 LDBL[142] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2793 LDBL[158] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2794 float1410 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2795 LDBL[190] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2796 LDBL[206] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2797 LDBL[222] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2798 LDBL[238] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2799 float1411 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=047e   word=15   wl=10 address=00af
m2800 float1412 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2801 LDBL[31] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2802 LDBL[47] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2803 LDBL[63] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2804 LDBL[79] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2805 LDBL[95] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2806 LDBL[111] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2807 float1413 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2808 float1414 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2809 float1415 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2810 LDBL[175] LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2811 float1416 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2812 float1417 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2813 float1418 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2814 float1419 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2815 float1420 LDWL[10] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f2a8   word=0   wl=11 address=00b0
m2816 float1421 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2817 float1422 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2818 float1423 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2819 LDBL[48] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2820 float1424 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2821 LDBL[80] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2822 float1425 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2823 LDBL[112] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2824 float1426 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2825 LDBL[144] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2826 float1427 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2827 float1428 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2828 LDBL[192] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2829 LDBL[208] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2830 LDBL[224] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2831 LDBL[240] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1a27   word=1   wl=11 address=00b1
m2832 LDBL[1] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2833 LDBL[17] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2834 LDBL[33] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2835 float1429 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2836 float1430 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2837 LDBL[81] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2838 float1431 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2839 float1432 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2840 float1433 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2841 LDBL[145] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2842 float1434 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2843 LDBL[177] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2844 LDBL[193] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2845 float1435 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2846 float1436 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2847 float1437 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0668   word=2   wl=11 address=00b2
m2848 float1438 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2849 float1439 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2850 float1440 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2851 LDBL[50] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2852 float1441 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2853 LDBL[82] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2854 LDBL[98] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2855 float1442 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2856 float1443 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2857 LDBL[146] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2858 LDBL[162] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2859 float1444 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2860 float1445 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2861 float1446 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2862 float1447 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2863 float1448 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8fff   word=3   wl=11 address=00b3
m2864 LDBL[3] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2865 LDBL[19] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2866 LDBL[35] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2867 LDBL[51] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2868 LDBL[67] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2869 LDBL[83] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2870 LDBL[99] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2871 LDBL[115] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2872 LDBL[131] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2873 LDBL[147] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2874 LDBL[163] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2875 LDBL[179] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2876 float1449 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2877 float1450 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2878 float1451 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2879 LDBL[243] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3a5c   word=4   wl=11 address=00b4
m2880 float1452 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2881 float1453 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2882 LDBL[36] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2883 LDBL[52] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2884 LDBL[68] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2885 float1454 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2886 LDBL[100] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2887 float1455 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2888 float1456 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2889 LDBL[148] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2890 float1457 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2891 LDBL[180] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2892 LDBL[196] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2893 LDBL[212] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2894 float1458 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2895 float1459 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7b14   word=5   wl=11 address=00b5
m2896 float1460 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2897 float1461 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2898 LDBL[37] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2899 float1462 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2900 LDBL[69] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2901 float1463 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2902 float1464 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2903 float1465 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2904 LDBL[133] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2905 LDBL[149] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2906 float1466 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2907 LDBL[181] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2908 LDBL[197] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2909 LDBL[213] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2910 LDBL[229] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2911 float1467 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=56f6   word=6   wl=11 address=00b6
m2912 float1468 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2913 LDBL[22] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2914 LDBL[38] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2915 float1469 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2916 LDBL[70] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2917 LDBL[86] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2918 LDBL[102] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2919 LDBL[118] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2920 float1470 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2921 LDBL[150] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2922 LDBL[166] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2923 float1471 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2924 LDBL[198] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2925 float1472 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2926 LDBL[230] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2927 float1473 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e350   word=7   wl=11 address=00b7
m2928 float1474 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2929 float1475 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2930 float1476 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2931 float1477 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2932 LDBL[71] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2933 float1478 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2934 LDBL[103] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2935 float1479 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2936 LDBL[135] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2937 LDBL[151] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2938 float1480 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2939 float1481 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2940 float1482 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2941 LDBL[215] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2942 LDBL[231] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2943 LDBL[247] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c02b   word=8   wl=11 address=00b8
m2944 LDBL[8] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2945 LDBL[24] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2946 float1483 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2947 LDBL[56] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2948 float1484 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2949 LDBL[88] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2950 float1485 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2951 float1486 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2952 float1487 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2953 float1488 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2954 float1489 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2955 float1490 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2956 float1491 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2957 float1492 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2958 LDBL[232] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2959 LDBL[248] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9f02   word=9   wl=11 address=00b9
m2960 float1493 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2961 LDBL[25] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2962 float1494 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2963 float1495 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2964 float1496 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2965 float1497 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2966 float1498 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2967 float1499 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2968 LDBL[137] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2969 LDBL[153] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2970 LDBL[169] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2971 LDBL[185] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2972 LDBL[201] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2973 float1500 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2974 float1501 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2975 LDBL[249] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=81fe   word=10   wl=11 address=00ba
m2976 float1502 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2977 LDBL[26] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2978 LDBL[42] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2979 LDBL[58] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2980 LDBL[74] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2981 LDBL[90] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2982 LDBL[106] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2983 LDBL[122] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2984 LDBL[138] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2985 float1503 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2986 float1504 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2987 float1505 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2988 float1506 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2989 float1507 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2990 float1508 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2991 LDBL[250] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f6df   word=11   wl=11 address=00bb
m2992 LDBL[11] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2993 LDBL[27] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2994 LDBL[43] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2995 LDBL[59] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2996 LDBL[75] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2997 float1509 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2998 LDBL[107] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m2999 LDBL[123] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3000 float1510 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3001 LDBL[155] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3002 LDBL[171] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3003 float1511 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3004 LDBL[203] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3005 LDBL[219] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3006 LDBL[235] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3007 LDBL[251] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=88cb   word=12   wl=11 address=00bc
m3008 LDBL[12] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3009 LDBL[28] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3010 float1512 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3011 LDBL[60] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3012 float1513 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3013 float1514 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3014 LDBL[108] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3015 LDBL[124] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3016 float1515 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3017 float1516 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3018 float1517 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3019 LDBL[188] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3020 float1518 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3021 float1519 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3022 float1520 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3023 LDBL[252] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=87c6   word=13   wl=11 address=00bd
m3024 float1521 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3025 LDBL[29] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3026 LDBL[45] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3027 float1522 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3028 float1523 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3029 float1524 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3030 LDBL[109] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3031 LDBL[125] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3032 LDBL[141] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3033 LDBL[157] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3034 LDBL[173] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3035 float1525 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3036 float1526 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3037 float1527 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3038 float1528 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3039 LDBL[253] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=39ff   word=14   wl=11 address=00be
m3040 LDBL[14] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3041 LDBL[30] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3042 LDBL[46] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3043 LDBL[62] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3044 LDBL[78] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3045 LDBL[94] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3046 LDBL[110] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3047 LDBL[126] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3048 LDBL[142] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3049 float1529 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3050 float1530 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3051 LDBL[190] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3052 LDBL[206] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3053 LDBL[222] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3054 float1531 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3055 float1532 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=879e   word=15   wl=11 address=00bf
m3056 float1533 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3057 LDBL[31] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3058 LDBL[47] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3059 LDBL[63] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3060 LDBL[79] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3061 float1534 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3062 float1535 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3063 LDBL[127] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3064 LDBL[143] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3065 LDBL[159] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3066 LDBL[175] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3067 float1536 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3068 float1537 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3069 float1538 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3070 float1539 LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3071 LDBL[255] LDWL[11] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b75e   word=0   wl=12 address=00c0
m3072 float1540 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3073 LDBL[16] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3074 LDBL[32] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3075 LDBL[48] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3076 LDBL[64] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3077 float1541 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3078 LDBL[96] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3079 float1542 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3080 LDBL[128] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3081 LDBL[144] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3082 LDBL[160] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3083 float1543 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3084 LDBL[192] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3085 LDBL[208] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3086 float1544 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3087 LDBL[240] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9f30   word=1   wl=12 address=00c1
m3088 float1545 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3089 float1546 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3090 float1547 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3091 float1548 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3092 LDBL[65] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3093 LDBL[81] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3094 float1549 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3095 float1550 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3096 LDBL[129] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3097 LDBL[145] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3098 LDBL[161] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3099 LDBL[177] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3100 LDBL[193] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3101 float1551 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3102 float1552 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3103 LDBL[241] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4de1   word=2   wl=12 address=00c2
m3104 LDBL[2] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3105 float1553 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3106 float1554 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3107 float1555 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3108 float1556 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3109 LDBL[82] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3110 LDBL[98] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3111 LDBL[114] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3112 LDBL[130] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3113 float1557 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3114 LDBL[162] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3115 LDBL[178] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3116 float1558 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3117 float1559 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3118 LDBL[226] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3119 float1560 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4bec   word=3   wl=12 address=00c3
m3120 float1561 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3121 float1562 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3122 LDBL[35] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3123 LDBL[51] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3124 float1563 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3125 LDBL[83] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3126 LDBL[99] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3127 LDBL[115] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3128 LDBL[131] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3129 LDBL[147] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3130 float1564 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3131 LDBL[179] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3132 float1565 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3133 float1566 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3134 LDBL[227] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3135 float1567 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=da53   word=4   wl=12 address=00c4
m3136 LDBL[4] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3137 LDBL[20] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3138 float1568 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3139 float1569 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3140 LDBL[68] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3141 float1570 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3142 LDBL[100] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3143 float1571 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3144 float1572 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3145 LDBL[148] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3146 float1573 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3147 LDBL[180] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3148 LDBL[196] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3149 float1574 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3150 LDBL[228] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3151 LDBL[244] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ef35   word=5   wl=12 address=00c5
m3152 LDBL[5] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3153 float1575 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3154 LDBL[37] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3155 float1576 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3156 LDBL[69] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3157 LDBL[85] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3158 float1577 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3159 float1578 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3160 LDBL[133] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3161 LDBL[149] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3162 LDBL[165] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3163 LDBL[181] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3164 float1579 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3165 LDBL[213] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3166 LDBL[229] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3167 LDBL[245] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=cafc   word=6   wl=12 address=00c6
m3168 float1580 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3169 float1581 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3170 LDBL[38] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3171 LDBL[54] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3172 LDBL[70] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3173 LDBL[86] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3174 LDBL[102] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3175 LDBL[118] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3176 float1582 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3177 LDBL[150] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3178 float1583 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3179 LDBL[182] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3180 float1584 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3181 float1585 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3182 LDBL[230] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3183 LDBL[246] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f3c5   word=7   wl=12 address=00c7
m3184 LDBL[7] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3185 float1586 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3186 LDBL[39] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3187 float1587 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3188 float1588 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3189 float1589 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3190 LDBL[103] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3191 LDBL[119] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3192 LDBL[135] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3193 LDBL[151] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3194 float1590 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3195 float1591 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3196 LDBL[199] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3197 LDBL[215] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3198 LDBL[231] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3199 LDBL[247] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0e24   word=8   wl=12 address=00c8
m3200 float1592 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3201 float1593 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3202 LDBL[40] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3203 float1594 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3204 float1595 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3205 LDBL[88] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3206 float1596 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3207 float1597 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3208 float1598 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3209 LDBL[152] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3210 LDBL[168] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3211 LDBL[184] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3212 float1599 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3213 float1600 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3214 float1601 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3215 float1602 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9c90   word=9   wl=12 address=00c9
m3216 float1603 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3217 float1604 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3218 float1605 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3219 float1606 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3220 LDBL[73] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3221 float1607 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3222 float1608 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3223 LDBL[121] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3224 float1609 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3225 float1610 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3226 LDBL[169] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3227 LDBL[185] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3228 LDBL[201] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3229 float1611 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3230 float1612 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3231 LDBL[249] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=415f   word=10   wl=12 address=00ca
m3232 LDBL[10] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3233 LDBL[26] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3234 LDBL[42] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3235 LDBL[58] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3236 LDBL[74] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3237 float1613 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3238 LDBL[106] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3239 float1614 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3240 LDBL[138] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3241 float1615 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3242 float1616 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3243 float1617 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3244 float1618 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3245 float1619 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3246 LDBL[234] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3247 float1620 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8c23   word=11   wl=12 address=00cb
m3248 LDBL[11] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3249 LDBL[27] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3250 float1621 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3251 float1622 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3252 float1623 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3253 LDBL[91] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3254 float1624 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3255 float1625 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3256 float1626 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3257 float1627 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3258 LDBL[171] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3259 LDBL[187] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3260 float1628 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3261 float1629 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3262 float1630 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3263 LDBL[251] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f57d   word=12   wl=12 address=00cc
m3264 LDBL[12] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3265 float1631 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3266 LDBL[44] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3267 LDBL[60] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3268 LDBL[76] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3269 LDBL[92] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3270 LDBL[108] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3271 float1632 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3272 LDBL[140] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3273 float1633 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3274 LDBL[172] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3275 float1634 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3276 LDBL[204] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3277 LDBL[220] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3278 LDBL[236] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3279 LDBL[252] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4281   word=13   wl=12 address=00cd
m3280 LDBL[13] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3281 float1635 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3282 float1636 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3283 float1637 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3284 float1638 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3285 float1639 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3286 float1640 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3287 LDBL[125] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3288 float1641 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3289 LDBL[157] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3290 float1642 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3291 float1643 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3292 float1644 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3293 float1645 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3294 LDBL[237] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3295 float1646 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ca01   word=14   wl=12 address=00ce
m3296 LDBL[14] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3297 float1647 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3298 float1648 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3299 float1649 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3300 float1650 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3301 float1651 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3302 float1652 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3303 float1653 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3304 float1654 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3305 LDBL[158] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3306 float1655 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3307 LDBL[190] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3308 float1656 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3309 float1657 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3310 LDBL[238] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3311 LDBL[254] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8662   word=15   wl=12 address=00cf
m3312 float1658 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3313 LDBL[31] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3314 float1659 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3315 float1660 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3316 float1661 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3317 LDBL[95] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3318 LDBL[111] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3319 float1662 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3320 float1663 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3321 LDBL[159] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3322 LDBL[175] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3323 float1664 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3324 float1665 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3325 float1666 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3326 float1667 LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3327 LDBL[255] LDWL[12] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2a1f   word=0   wl=13 address=00d0
m3328 LDBL[0] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3329 LDBL[16] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3330 LDBL[32] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3331 LDBL[48] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3332 LDBL[64] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3333 float1668 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3334 float1669 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3335 float1670 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3336 float1671 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3337 LDBL[144] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3338 float1672 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3339 LDBL[176] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3340 float1673 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3341 LDBL[208] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3342 float1674 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3343 float1675 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=035d   word=1   wl=13 address=00d1
m3344 LDBL[1] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3345 float1676 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3346 LDBL[33] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3347 LDBL[49] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3348 LDBL[65] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3349 float1677 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3350 LDBL[97] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3351 float1678 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3352 LDBL[129] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3353 LDBL[145] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3354 float1679 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3355 float1680 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3356 float1681 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3357 float1682 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3358 float1683 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3359 float1684 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fd1f   word=2   wl=13 address=00d2
m3360 LDBL[2] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3361 LDBL[18] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3362 LDBL[34] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3363 LDBL[50] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3364 LDBL[66] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3365 float1685 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3366 float1686 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3367 float1687 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3368 LDBL[130] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3369 float1688 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3370 LDBL[162] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3371 LDBL[178] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3372 LDBL[194] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3373 LDBL[210] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3374 LDBL[226] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3375 LDBL[242] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=045a   word=3   wl=13 address=00d3
m3376 float1689 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3377 LDBL[19] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3378 float1690 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3379 LDBL[51] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3380 LDBL[67] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3381 float1691 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3382 LDBL[99] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3383 float1692 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3384 float1693 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3385 float1694 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3386 LDBL[163] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3387 float1695 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3388 float1696 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3389 float1697 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3390 float1698 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3391 float1699 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9980   word=4   wl=13 address=00d4
m3392 float1700 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3393 float1701 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3394 float1702 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3395 float1703 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3396 float1704 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3397 float1705 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3398 float1706 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3399 LDBL[116] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3400 LDBL[132] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3401 float1707 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3402 float1708 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3403 LDBL[180] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3404 LDBL[196] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3405 float1709 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3406 float1710 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3407 LDBL[244] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a7a2   word=5   wl=13 address=00d5
m3408 float1711 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3409 LDBL[21] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3410 float1712 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3411 float1713 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3412 float1714 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3413 LDBL[85] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3414 float1715 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3415 LDBL[117] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3416 LDBL[133] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3417 LDBL[149] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3418 LDBL[165] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3419 float1716 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3420 float1717 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3421 LDBL[213] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3422 float1718 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3423 LDBL[245] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=230c   word=6   wl=13 address=00d6
m3424 float1719 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3425 float1720 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3426 LDBL[38] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3427 LDBL[54] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3428 float1721 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3429 float1722 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3430 float1723 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3431 float1724 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3432 LDBL[134] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3433 LDBL[150] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3434 float1725 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3435 float1726 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3436 float1727 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3437 LDBL[214] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3438 float1728 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3439 float1729 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=bc03   word=7   wl=13 address=00d7
m3440 LDBL[7] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3441 LDBL[23] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3442 float1730 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3443 float1731 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3444 float1732 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3445 float1733 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3446 float1734 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3447 float1735 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3448 float1736 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3449 float1737 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3450 LDBL[167] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3451 LDBL[183] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3452 LDBL[199] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3453 LDBL[215] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3454 float1738 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3455 LDBL[247] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3dbd   word=8   wl=13 address=00d8
m3456 LDBL[8] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3457 float1739 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3458 LDBL[40] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3459 LDBL[56] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3460 LDBL[72] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3461 LDBL[88] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3462 float1740 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3463 LDBL[120] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3464 LDBL[136] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3465 float1741 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3466 LDBL[168] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3467 LDBL[184] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3468 LDBL[200] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3469 LDBL[216] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3470 float1742 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3471 float1743 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ad0f   word=9   wl=13 address=00d9
m3472 LDBL[9] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3473 LDBL[25] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3474 LDBL[41] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3475 LDBL[57] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3476 float1744 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3477 float1745 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3478 float1746 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3479 float1747 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3480 LDBL[137] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3481 float1748 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3482 LDBL[169] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3483 LDBL[185] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3484 float1749 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3485 LDBL[217] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3486 float1750 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3487 LDBL[249] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=39df   word=10   wl=13 address=00da
m3488 LDBL[10] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3489 LDBL[26] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3490 LDBL[42] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3491 LDBL[58] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3492 LDBL[74] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3493 float1751 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3494 LDBL[106] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3495 LDBL[122] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3496 LDBL[138] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3497 float1752 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3498 float1753 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3499 LDBL[186] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3500 LDBL[202] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3501 LDBL[218] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3502 float1754 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3503 float1755 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=22a1   word=11   wl=13 address=00db
m3504 LDBL[11] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3505 float1756 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3506 float1757 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3507 float1758 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3508 float1759 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3509 LDBL[91] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3510 float1760 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3511 LDBL[123] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3512 float1761 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3513 LDBL[155] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3514 float1762 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3515 float1763 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3516 float1764 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3517 LDBL[219] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3518 float1765 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3519 float1766 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6cca   word=12   wl=13 address=00dc
m3520 float1767 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3521 LDBL[28] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3522 float1768 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3523 LDBL[60] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3524 float1769 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3525 float1770 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3526 LDBL[108] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3527 LDBL[124] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3528 float1771 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3529 float1772 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3530 LDBL[172] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3531 LDBL[188] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3532 float1773 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3533 LDBL[220] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3534 LDBL[236] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3535 float1774 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c1c9   word=13   wl=13 address=00dd
m3536 LDBL[13] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3537 float1775 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3538 float1776 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3539 LDBL[61] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3540 float1777 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3541 float1778 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3542 LDBL[109] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3543 LDBL[125] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3544 LDBL[141] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3545 float1779 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3546 float1780 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3547 float1781 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3548 float1782 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3549 float1783 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3550 LDBL[237] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3551 LDBL[253] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a1a9   word=14   wl=13 address=00de
m3552 LDBL[14] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3553 float1784 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3554 float1785 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3555 LDBL[62] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3556 float1786 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3557 LDBL[94] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3558 float1787 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3559 LDBL[126] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3560 LDBL[142] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3561 float1788 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3562 float1789 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3563 float1790 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3564 float1791 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3565 LDBL[222] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3566 float1792 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3567 LDBL[254] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6607   word=15   wl=13 address=00df
m3568 LDBL[15] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3569 LDBL[31] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3570 LDBL[47] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3571 float1793 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3572 float1794 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3573 float1795 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3574 float1796 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3575 float1797 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3576 float1798 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3577 LDBL[159] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3578 LDBL[175] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3579 float1799 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3580 float1800 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3581 LDBL[223] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3582 LDBL[239] LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3583 float1801 LDWL[13] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d846   word=0   wl=14 address=00e0
m3584 float1802 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3585 LDBL[16] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3586 LDBL[32] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3587 float1803 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3588 float1804 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3589 float1805 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3590 LDBL[96] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3591 float1806 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3592 float1807 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3593 float1808 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3594 float1809 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3595 LDBL[176] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3596 LDBL[192] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3597 float1810 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3598 LDBL[224] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3599 LDBL[240] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5c5d   word=1   wl=14 address=00e1
m3600 LDBL[1] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3601 float1811 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3602 LDBL[33] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3603 LDBL[49] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3604 LDBL[65] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3605 float1812 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3606 LDBL[97] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3607 float1813 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3608 float1814 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3609 float1815 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3610 LDBL[161] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3611 LDBL[177] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3612 LDBL[193] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3613 float1816 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3614 LDBL[225] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3615 float1817 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=acca   word=2   wl=14 address=00e2
m3616 float1818 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3617 LDBL[18] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3618 float1819 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3619 LDBL[50] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3620 float1820 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3621 float1821 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3622 LDBL[98] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3623 LDBL[114] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3624 float1822 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3625 float1823 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3626 LDBL[162] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3627 LDBL[178] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3628 float1824 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3629 LDBL[210] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3630 float1825 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3631 LDBL[242] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=357f   word=3   wl=14 address=00e3
m3632 LDBL[3] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3633 LDBL[19] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3634 LDBL[35] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3635 LDBL[51] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3636 LDBL[67] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3637 LDBL[83] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3638 LDBL[99] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3639 float1826 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3640 LDBL[131] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3641 float1827 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3642 LDBL[163] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3643 float1828 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3644 LDBL[195] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3645 LDBL[211] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3646 float1829 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3647 float1830 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b1a4   word=4   wl=14 address=00e4
m3648 float1831 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3649 float1832 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3650 LDBL[36] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3651 float1833 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3652 float1834 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3653 LDBL[84] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3654 float1835 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3655 LDBL[116] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3656 LDBL[132] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3657 float1836 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3658 float1837 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3659 float1838 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3660 LDBL[196] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3661 LDBL[212] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3662 float1839 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3663 LDBL[244] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=bbd7   word=5   wl=14 address=00e5
m3664 LDBL[5] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3665 LDBL[21] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3666 LDBL[37] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3667 float1840 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3668 LDBL[69] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3669 float1841 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3670 LDBL[101] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3671 LDBL[117] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3672 LDBL[133] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3673 LDBL[149] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3674 float1842 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3675 LDBL[181] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3676 LDBL[197] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3677 LDBL[213] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3678 float1843 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3679 LDBL[245] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4082   word=6   wl=14 address=00e6
m3680 float1844 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3681 LDBL[22] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3682 float1845 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3683 float1846 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3684 float1847 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3685 float1848 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3686 float1849 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3687 LDBL[118] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3688 float1850 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3689 float1851 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3690 float1852 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3691 float1853 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3692 float1854 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3693 float1855 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3694 LDBL[230] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3695 float1856 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5bcf   word=7   wl=14 address=00e7
m3696 LDBL[7] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3697 LDBL[23] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3698 LDBL[39] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3699 LDBL[55] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3700 float1857 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3701 float1858 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3702 LDBL[103] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3703 LDBL[119] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3704 LDBL[135] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3705 LDBL[151] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3706 float1859 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3707 LDBL[183] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3708 LDBL[199] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3709 float1860 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3710 LDBL[231] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3711 float1861 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2387   word=8   wl=14 address=00e8
m3712 LDBL[8] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3713 LDBL[24] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3714 LDBL[40] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3715 float1862 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3716 float1863 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3717 float1864 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3718 float1865 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3719 LDBL[120] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3720 LDBL[136] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3721 LDBL[152] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3722 float1866 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3723 float1867 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3724 float1868 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3725 LDBL[216] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3726 float1869 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3727 float1870 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d27a   word=9   wl=14 address=00e9
m3728 float1871 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3729 LDBL[25] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3730 float1872 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3731 LDBL[57] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3732 LDBL[73] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3733 LDBL[89] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3734 LDBL[105] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3735 float1873 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3736 float1874 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3737 LDBL[153] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3738 float1875 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3739 float1876 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3740 LDBL[201] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3741 float1877 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3742 LDBL[233] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3743 LDBL[249] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1fc8   word=10   wl=14 address=00ea
m3744 float1878 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3745 float1879 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3746 float1880 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3747 LDBL[58] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3748 float1881 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3749 float1882 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3750 LDBL[106] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3751 LDBL[122] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3752 LDBL[138] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3753 LDBL[154] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3754 LDBL[170] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3755 LDBL[186] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3756 LDBL[202] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3757 float1883 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3758 float1884 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3759 float1885 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=de69   word=11   wl=14 address=00eb
m3760 LDBL[11] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3761 float1886 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3762 float1887 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3763 LDBL[59] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3764 float1888 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3765 LDBL[91] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3766 LDBL[107] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3767 float1889 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3768 float1890 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3769 LDBL[155] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3770 LDBL[171] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3771 LDBL[187] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3772 LDBL[203] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3773 float1891 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3774 LDBL[235] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3775 LDBL[251] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8121   word=12   wl=14 address=00ec
m3776 LDBL[12] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3777 float1892 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3778 float1893 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3779 float1894 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3780 float1895 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3781 LDBL[92] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3782 float1896 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3783 float1897 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3784 LDBL[140] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3785 float1898 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3786 float1899 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3787 float1900 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3788 float1901 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3789 float1902 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3790 float1903 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3791 LDBL[252] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=190b   word=13   wl=14 address=00ed
m3792 LDBL[13] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3793 LDBL[29] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3794 float1904 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3795 LDBL[61] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3796 float1905 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3797 float1906 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3798 float1907 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3799 float1908 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3800 LDBL[141] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3801 float1909 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3802 float1910 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3803 LDBL[189] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3804 LDBL[205] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3805 float1911 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3806 float1912 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3807 float1913 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c1a0   word=14   wl=14 address=00ee
m3808 float1914 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3809 float1915 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3810 float1916 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3811 float1917 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3812 float1918 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3813 LDBL[94] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3814 float1919 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3815 LDBL[126] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3816 LDBL[142] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3817 float1920 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3818 float1921 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3819 float1922 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3820 float1923 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3821 float1924 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3822 LDBL[238] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3823 LDBL[254] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e8f8   word=15   wl=14 address=00ef
m3824 float1925 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3825 float1926 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3826 float1927 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3827 LDBL[63] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3828 LDBL[79] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3829 LDBL[95] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3830 LDBL[111] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3831 LDBL[127] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3832 float1928 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3833 float1929 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3834 float1930 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3835 LDBL[191] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3836 float1931 LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3837 LDBL[223] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3838 LDBL[239] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3839 LDBL[255] LDWL[14] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fa05   word=0   wl=15 address=00f0
m3840 LDBL[0] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3841 float1932 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3842 LDBL[32] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3843 float1933 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3844 float1934 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3845 float1935 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3846 float1936 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3847 float1937 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3848 float1938 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3849 LDBL[144] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3850 float1939 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3851 LDBL[176] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3852 LDBL[192] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3853 LDBL[208] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3854 LDBL[224] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3855 LDBL[240] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=43a7   word=1   wl=15 address=00f1
m3856 LDBL[1] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3857 LDBL[17] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3858 LDBL[33] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3859 float1940 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3860 float1941 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3861 LDBL[81] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3862 float1942 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3863 LDBL[113] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3864 LDBL[129] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3865 LDBL[145] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3866 float1943 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3867 float1944 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3868 float1945 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3869 float1946 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3870 LDBL[225] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3871 float1947 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c28f   word=2   wl=15 address=00f2
m3872 LDBL[2] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3873 LDBL[18] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3874 LDBL[34] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3875 LDBL[50] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3876 float1948 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3877 float1949 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3878 float1950 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3879 LDBL[114] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3880 float1951 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3881 LDBL[146] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3882 float1952 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3883 float1953 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3884 float1954 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3885 float1955 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3886 LDBL[226] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3887 LDBL[242] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9278   word=3   wl=15 address=00f3
m3888 float1956 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3889 float1957 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3890 float1958 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3891 LDBL[51] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3892 LDBL[67] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3893 LDBL[83] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3894 LDBL[99] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3895 float1959 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3896 float1960 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3897 LDBL[147] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3898 float1961 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3899 float1962 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3900 LDBL[195] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3901 float1963 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3902 float1964 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3903 LDBL[243] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=953c   word=4   wl=15 address=00f4
m3904 float1965 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3905 float1966 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3906 LDBL[36] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3907 LDBL[52] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3908 LDBL[68] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3909 LDBL[84] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3910 float1967 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3911 float1968 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3912 LDBL[132] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3913 float1969 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3914 LDBL[164] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3915 float1970 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3916 LDBL[196] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3917 float1971 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3918 float1972 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3919 LDBL[244] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b2d4   word=5   wl=15 address=00f5
m3920 float1973 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3921 float1974 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3922 LDBL[37] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3923 float1975 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3924 LDBL[69] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3925 float1976 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3926 LDBL[101] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3927 LDBL[117] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3928 float1977 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3929 LDBL[149] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3930 float1978 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3931 float1979 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3932 LDBL[197] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3933 LDBL[213] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3934 float1980 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3935 LDBL[245] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c108   word=6   wl=15 address=00f6
m3936 float1981 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3937 float1982 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3938 float1983 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3939 LDBL[54] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3940 float1984 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3941 float1985 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3942 float1986 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3943 float1987 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3944 LDBL[134] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3945 float1988 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3946 float1989 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3947 float1990 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3948 float1991 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3949 float1992 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3950 LDBL[230] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3951 LDBL[246] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f848   word=7   wl=15 address=00f7
m3952 float1993 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3953 float1994 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3954 float1995 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3955 LDBL[55] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3956 float1996 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3957 float1997 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3958 LDBL[103] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3959 float1998 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3960 float1999 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3961 float2000 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3962 float2001 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3963 LDBL[183] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3964 LDBL[199] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3965 LDBL[215] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3966 LDBL[231] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3967 LDBL[247] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f0ce   word=8   wl=15 address=00f8
m3968 float2002 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3969 LDBL[24] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3970 LDBL[40] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3971 LDBL[56] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3972 float2003 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3973 float2004 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3974 LDBL[104] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3975 LDBL[120] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3976 float2005 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3977 float2006 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3978 float2007 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3979 float2008 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3980 LDBL[200] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3981 LDBL[216] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3982 LDBL[232] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3983 LDBL[248] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6bf4   word=9   wl=15 address=00f9
m3984 float2009 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3985 float2010 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3986 LDBL[41] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3987 float2011 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3988 LDBL[73] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3989 LDBL[89] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3990 LDBL[105] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3991 LDBL[121] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3992 LDBL[137] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3993 LDBL[153] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3994 float2012 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3995 LDBL[185] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3996 float2013 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3997 LDBL[217] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3998 LDBL[233] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m3999 float2014 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e3d3   word=10   wl=15 address=00fa
m4000 LDBL[10] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4001 LDBL[26] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4002 float2015 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4003 float2016 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4004 LDBL[74] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4005 float2017 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4006 LDBL[106] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4007 LDBL[122] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4008 LDBL[138] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4009 LDBL[154] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4010 float2018 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4011 float2019 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4012 float2020 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4013 LDBL[218] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4014 LDBL[234] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4015 LDBL[250] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=592e   word=11   wl=15 address=00fb
m4016 float2021 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4017 LDBL[27] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4018 LDBL[43] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4019 LDBL[59] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4020 float2022 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4021 LDBL[91] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4022 float2023 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4023 float2024 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4024 LDBL[139] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4025 float2025 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4026 float2026 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4027 LDBL[187] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4028 LDBL[203] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4029 float2027 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4030 LDBL[235] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4031 float2028 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=269e   word=12   wl=15 address=00fc
m4032 float2029 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4033 LDBL[28] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4034 LDBL[44] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4035 LDBL[60] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4036 LDBL[76] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4037 float2030 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4038 float2031 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4039 LDBL[124] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4040 float2032 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4041 LDBL[156] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4042 LDBL[172] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4043 float2033 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4044 float2034 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4045 LDBL[220] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4046 float2035 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4047 float2036 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2db7   word=13   wl=15 address=00fd
m4048 LDBL[13] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4049 LDBL[29] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4050 LDBL[45] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4051 float2037 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4052 LDBL[77] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4053 LDBL[93] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4054 float2038 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4055 LDBL[125] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4056 LDBL[141] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4057 float2039 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4058 LDBL[173] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4059 LDBL[189] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4060 float2040 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4061 LDBL[221] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4062 float2041 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4063 float2042 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=dae2   word=14   wl=15 address=00fe
m4064 float2043 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4065 LDBL[30] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4066 float2044 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4067 float2045 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4068 float2046 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4069 LDBL[94] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4070 LDBL[110] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4071 LDBL[126] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4072 float2047 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4073 LDBL[158] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4074 float2048 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4075 LDBL[190] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4076 LDBL[206] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4077 float2049 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4078 LDBL[238] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4079 LDBL[254] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7076   word=15   wl=15 address=00ff
m4080 float2050 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4081 LDBL[31] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4082 LDBL[47] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4083 float2051 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4084 LDBL[79] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4085 LDBL[95] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4086 LDBL[111] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4087 float2052 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4088 float2053 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4089 float2054 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4090 float2055 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4091 float2056 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4092 LDBL[207] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4093 LDBL[223] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4094 LDBL[239] LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4095 float2057 LDWL[15] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=032f   word=0   wl=16 address=0100
m4096 LDBL[0] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4097 LDBL[16] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4098 LDBL[32] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4099 LDBL[48] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4100 float2058 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4101 LDBL[80] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4102 float2059 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4103 float2060 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4104 LDBL[128] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4105 LDBL[144] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4106 float2061 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4107 float2062 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4108 float2063 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4109 float2064 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4110 float2065 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4111 float2066 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=95ce   word=1   wl=16 address=0101
m4112 float2067 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4113 LDBL[17] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4114 LDBL[33] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4115 LDBL[49] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4116 float2068 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4117 float2069 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4118 LDBL[97] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4119 LDBL[113] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4120 LDBL[129] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4121 float2070 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4122 LDBL[161] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4123 float2071 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4124 LDBL[193] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4125 float2072 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4126 float2073 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4127 LDBL[241] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1855   word=2   wl=16 address=0102
m4128 LDBL[2] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4129 float2074 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4130 LDBL[34] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4131 float2075 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4132 LDBL[66] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4133 float2076 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4134 LDBL[98] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4135 float2077 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4136 float2078 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4137 float2079 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4138 float2080 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4139 LDBL[178] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4140 LDBL[194] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4141 float2081 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4142 float2082 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4143 float2083 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0d17   word=3   wl=16 address=0103
m4144 LDBL[3] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4145 LDBL[19] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4146 LDBL[35] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4147 float2084 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4148 LDBL[67] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4149 float2085 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4150 float2086 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4151 float2087 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4152 LDBL[131] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4153 float2088 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4154 LDBL[163] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4155 LDBL[179] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4156 float2089 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4157 float2090 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4158 float2091 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4159 float2092 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ed6d   word=4   wl=16 address=0104
m4160 LDBL[4] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4161 float2093 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4162 LDBL[36] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4163 LDBL[52] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4164 float2094 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4165 LDBL[84] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4166 LDBL[100] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4167 float2095 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4168 LDBL[132] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4169 float2096 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4170 LDBL[164] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4171 LDBL[180] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4172 float2097 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4173 LDBL[212] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4174 LDBL[228] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4175 LDBL[244] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1207   word=5   wl=16 address=0105
m4176 LDBL[5] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4177 LDBL[21] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4178 LDBL[37] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4179 float2098 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4180 float2099 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4181 float2100 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4182 float2101 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4183 float2102 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4184 float2103 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4185 LDBL[149] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4186 float2104 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4187 float2105 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4188 LDBL[197] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4189 float2106 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4190 float2107 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4191 float2108 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5147   word=6   wl=16 address=0106
m4192 LDBL[6] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4193 LDBL[22] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4194 LDBL[38] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4195 float2109 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4196 float2110 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4197 float2111 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4198 LDBL[102] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4199 float2112 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4200 LDBL[134] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4201 float2113 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4202 float2114 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4203 float2115 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4204 LDBL[198] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4205 float2116 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4206 LDBL[230] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4207 float2117 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2717   word=7   wl=16 address=0107
m4208 LDBL[7] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4209 LDBL[23] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4210 LDBL[39] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4211 float2118 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4212 LDBL[71] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4213 float2119 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4214 float2120 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4215 float2121 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4216 LDBL[135] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4217 LDBL[151] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4218 LDBL[167] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4219 float2122 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4220 float2123 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4221 LDBL[215] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4222 float2124 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4223 float2125 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7fbd   word=8   wl=16 address=0108
m4224 LDBL[8] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4225 float2126 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4226 LDBL[40] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4227 LDBL[56] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4228 LDBL[72] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4229 LDBL[88] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4230 float2127 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4231 LDBL[120] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4232 LDBL[136] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4233 LDBL[152] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4234 LDBL[168] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4235 LDBL[184] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4236 LDBL[200] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4237 LDBL[216] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4238 LDBL[232] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4239 float2128 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2ccf   word=9   wl=16 address=0109
m4240 LDBL[9] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4241 LDBL[25] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4242 LDBL[41] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4243 LDBL[57] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4244 float2129 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4245 float2130 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4246 LDBL[105] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4247 LDBL[121] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4248 float2131 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4249 float2132 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4250 LDBL[169] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4251 LDBL[185] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4252 float2133 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4253 LDBL[217] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4254 float2134 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4255 float2135 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=51a8   word=10   wl=16 address=010a
m4256 float2136 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4257 float2137 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4258 float2138 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4259 LDBL[58] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4260 float2139 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4261 LDBL[90] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4262 float2140 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4263 LDBL[122] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4264 LDBL[138] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4265 float2141 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4266 float2142 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4267 float2143 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4268 LDBL[202] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4269 float2144 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4270 LDBL[234] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4271 float2145 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5bfe   word=11   wl=16 address=010b
m4272 float2146 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4273 LDBL[27] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4274 LDBL[43] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4275 LDBL[59] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4276 LDBL[75] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4277 LDBL[91] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4278 LDBL[107] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4279 LDBL[123] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4280 LDBL[139] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4281 LDBL[155] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4282 float2147 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4283 LDBL[187] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4284 LDBL[203] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4285 float2148 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4286 LDBL[235] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4287 float2149 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9509   word=12   wl=16 address=010c
m4288 LDBL[12] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4289 float2150 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4290 float2151 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4291 LDBL[60] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4292 float2152 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4293 float2153 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4294 float2154 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4295 float2155 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4296 LDBL[140] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4297 float2156 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4298 LDBL[172] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4299 float2157 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4300 LDBL[204] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4301 float2158 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4302 float2159 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4303 LDBL[252] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2321   word=13   wl=16 address=010d
m4304 LDBL[13] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4305 float2160 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4306 float2161 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4307 float2162 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4308 float2163 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4309 LDBL[93] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4310 float2164 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4311 float2165 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4312 LDBL[141] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4313 LDBL[157] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4314 float2166 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4315 float2167 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4316 float2168 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4317 LDBL[221] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4318 float2169 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4319 float2170 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3454   word=14   wl=16 address=010e
m4320 float2171 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4321 float2172 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4322 LDBL[46] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4323 float2173 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4324 LDBL[78] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4325 float2174 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4326 LDBL[110] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4327 float2175 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4328 float2176 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4329 float2177 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4330 LDBL[174] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4331 float2178 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4332 LDBL[206] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4333 LDBL[222] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4334 float2179 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4335 float2180 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ca87   word=15   wl=16 address=010f
m4336 LDBL[15] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4337 LDBL[31] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4338 LDBL[47] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4339 float2181 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4340 float2182 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4341 float2183 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4342 float2184 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4343 LDBL[127] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4344 float2185 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4345 LDBL[159] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4346 float2186 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4347 LDBL[191] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4348 float2187 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4349 float2188 LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4350 LDBL[239] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4351 LDBL[255] LDWL[16] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=da17   word=0   wl=17 address=0110
m4352 LDBL[0] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4353 LDBL[16] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4354 LDBL[32] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4355 float2189 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4356 LDBL[64] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4357 float2190 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4358 float2191 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4359 float2192 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4360 float2193 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4361 LDBL[144] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4362 float2194 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4363 LDBL[176] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4364 LDBL[192] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4365 float2195 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4366 LDBL[224] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4367 LDBL[240] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7404   word=1   wl=17 address=0111
m4368 float2196 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4369 float2197 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4370 LDBL[33] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4371 float2198 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4372 float2199 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4373 float2200 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4374 float2201 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4375 float2202 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4376 float2203 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4377 float2204 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4378 LDBL[161] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4379 float2205 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4380 LDBL[193] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4381 LDBL[209] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4382 LDBL[225] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4383 float2206 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=32bc   word=2   wl=17 address=0112
m4384 float2207 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4385 float2208 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4386 LDBL[34] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4387 LDBL[50] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4388 LDBL[66] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4389 LDBL[82] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4390 float2209 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4391 LDBL[114] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4392 float2210 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4393 LDBL[146] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4394 float2211 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4395 float2212 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4396 LDBL[194] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4397 LDBL[210] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4398 float2213 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4399 float2214 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a32a   word=3   wl=17 address=0113
m4400 float2215 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4401 LDBL[19] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4402 float2216 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4403 LDBL[51] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4404 float2217 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4405 LDBL[83] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4406 float2218 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4407 float2219 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4408 LDBL[131] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4409 LDBL[147] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4410 float2220 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4411 float2221 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4412 float2222 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4413 LDBL[211] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4414 float2223 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4415 LDBL[243] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e6a6   word=4   wl=17 address=0114
m4416 float2224 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4417 LDBL[20] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4418 LDBL[36] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4419 float2225 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4420 float2226 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4421 LDBL[84] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4422 float2227 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4423 LDBL[116] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4424 float2228 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4425 LDBL[148] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4426 LDBL[164] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4427 float2229 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4428 float2230 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4429 LDBL[212] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4430 LDBL[228] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4431 LDBL[244] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5392   word=5   wl=17 address=0115
m4432 float2231 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4433 LDBL[21] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4434 float2232 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4435 float2233 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4436 LDBL[69] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4437 float2234 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4438 float2235 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4439 LDBL[117] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4440 LDBL[133] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4441 LDBL[149] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4442 float2236 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4443 float2237 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4444 LDBL[197] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4445 float2238 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4446 LDBL[229] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4447 float2239 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7340   word=6   wl=17 address=0116
m4448 float2240 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4449 float2241 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4450 float2242 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4451 float2243 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4452 float2244 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4453 float2245 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4454 LDBL[102] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4455 float2246 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4456 LDBL[134] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4457 LDBL[150] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4458 float2247 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4459 float2248 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4460 LDBL[198] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4461 LDBL[214] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4462 LDBL[230] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4463 float2249 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8e0f   word=7   wl=17 address=0117
m4464 LDBL[7] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4465 LDBL[23] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4466 LDBL[39] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4467 LDBL[55] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4468 float2250 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4469 float2251 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4470 float2252 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4471 float2253 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4472 float2254 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4473 LDBL[151] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4474 LDBL[167] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4475 LDBL[183] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4476 float2255 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4477 float2256 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4478 float2257 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4479 LDBL[247] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=02f4   word=8   wl=17 address=0118
m4480 float2258 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4481 float2259 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4482 LDBL[40] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4483 float2260 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4484 LDBL[72] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4485 LDBL[88] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4486 LDBL[104] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4487 LDBL[120] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4488 float2261 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4489 LDBL[152] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4490 float2262 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4491 float2263 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4492 float2264 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4493 float2265 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4494 float2266 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4495 float2267 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=bba5   word=9   wl=17 address=0119
m4496 LDBL[9] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4497 float2268 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4498 LDBL[41] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4499 float2269 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4500 float2270 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4501 LDBL[89] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4502 float2271 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4503 LDBL[121] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4504 LDBL[137] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4505 LDBL[153] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4506 float2272 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4507 LDBL[185] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4508 LDBL[201] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4509 LDBL[217] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4510 float2273 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4511 LDBL[249] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e788   word=10   wl=17 address=011a
m4512 float2274 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4513 float2275 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4514 float2276 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4515 LDBL[58] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4516 float2277 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4517 float2278 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4518 float2279 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4519 LDBL[122] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4520 LDBL[138] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4521 LDBL[154] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4522 LDBL[170] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4523 float2280 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4524 float2281 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4525 LDBL[218] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4526 LDBL[234] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4527 LDBL[250] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2bdd   word=11   wl=17 address=011b
m4528 LDBL[11] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4529 float2282 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4530 LDBL[43] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4531 LDBL[59] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4532 LDBL[75] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4533 float2283 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4534 LDBL[107] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4535 LDBL[123] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4536 LDBL[139] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4537 LDBL[155] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4538 float2284 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4539 LDBL[187] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4540 float2285 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4541 LDBL[219] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4542 float2286 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4543 float2287 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=acfd   word=12   wl=17 address=011c
m4544 LDBL[12] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4545 float2288 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4546 LDBL[44] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4547 LDBL[60] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4548 LDBL[76] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4549 LDBL[92] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4550 LDBL[108] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4551 LDBL[124] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4552 float2289 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4553 float2290 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4554 LDBL[172] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4555 LDBL[188] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4556 float2291 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4557 LDBL[220] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4558 float2292 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4559 LDBL[252] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0986   word=13   wl=17 address=011d
m4560 float2293 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4561 LDBL[29] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4562 LDBL[45] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4563 float2294 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4564 float2295 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4565 float2296 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4566 float2297 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4567 LDBL[125] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4568 LDBL[141] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4569 float2298 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4570 float2299 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4571 LDBL[189] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4572 float2300 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4573 float2301 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4574 float2302 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4575 float2303 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=30bd   word=14   wl=17 address=011e
m4576 LDBL[14] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4577 float2304 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4578 LDBL[46] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4579 LDBL[62] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4580 LDBL[78] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4581 LDBL[94] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4582 float2305 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4583 LDBL[126] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4584 float2306 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4585 float2307 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4586 float2308 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4587 float2309 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4588 LDBL[206] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4589 LDBL[222] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4590 float2310 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4591 float2311 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=24e2   word=15   wl=17 address=011f
m4592 float2312 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4593 LDBL[31] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4594 float2313 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4595 float2314 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4596 float2315 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4597 LDBL[95] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4598 LDBL[111] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4599 LDBL[127] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4600 float2316 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4601 float2317 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4602 LDBL[175] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4603 float2318 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4604 float2319 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4605 LDBL[223] LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4606 float2320 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4607 float2321 LDWL[17] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c129   word=0   wl=18 address=0120
m4608 LDBL[0] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4609 float2322 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4610 float2323 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4611 LDBL[48] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4612 float2324 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4613 LDBL[80] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4614 float2325 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4615 float2326 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4616 LDBL[128] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4617 float2327 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4618 float2328 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4619 float2329 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4620 float2330 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4621 float2331 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4622 LDBL[224] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4623 LDBL[240] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e8de   word=1   wl=18 address=0121
m4624 float2332 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4625 LDBL[17] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4626 LDBL[33] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4627 LDBL[49] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4628 LDBL[65] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4629 float2333 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4630 LDBL[97] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4631 LDBL[113] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4632 float2334 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4633 float2335 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4634 float2336 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4635 LDBL[177] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4636 float2337 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4637 LDBL[209] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4638 LDBL[225] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4639 LDBL[241] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=dfe7   word=2   wl=18 address=0122
m4640 LDBL[2] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4641 LDBL[18] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4642 LDBL[34] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4643 float2338 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4644 float2339 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4645 LDBL[82] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4646 LDBL[98] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4647 LDBL[114] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4648 LDBL[130] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4649 LDBL[146] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4650 LDBL[162] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4651 LDBL[178] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4652 LDBL[194] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4653 float2340 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4654 LDBL[226] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4655 LDBL[242] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5f4a   word=3   wl=18 address=0123
m4656 float2341 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4657 LDBL[19] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4658 float2342 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4659 LDBL[51] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4660 float2343 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4661 float2344 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4662 LDBL[99] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4663 float2345 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4664 LDBL[131] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4665 LDBL[147] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4666 LDBL[163] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4667 LDBL[179] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4668 LDBL[195] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4669 float2346 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4670 LDBL[227] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4671 float2347 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=177e   word=4   wl=18 address=0124
m4672 float2348 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4673 LDBL[20] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4674 LDBL[36] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4675 LDBL[52] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4676 LDBL[68] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4677 LDBL[84] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4678 LDBL[100] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4679 float2349 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4680 LDBL[132] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4681 LDBL[148] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4682 LDBL[164] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4683 float2350 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4684 LDBL[196] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4685 float2351 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4686 float2352 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4687 float2353 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=37bc   word=5   wl=18 address=0125
m4688 float2354 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4689 float2355 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4690 LDBL[37] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4691 LDBL[53] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4692 LDBL[69] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4693 LDBL[85] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4694 float2356 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4695 LDBL[117] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4696 LDBL[133] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4697 LDBL[149] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4698 LDBL[165] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4699 float2357 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4700 LDBL[197] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4701 LDBL[213] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4702 float2358 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4703 float2359 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=99c2   word=6   wl=18 address=0126
m4704 float2360 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4705 LDBL[22] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4706 float2361 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4707 float2362 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4708 float2363 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4709 float2364 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4710 LDBL[102] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4711 LDBL[118] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4712 LDBL[134] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4713 float2365 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4714 float2366 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4715 LDBL[182] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4716 LDBL[198] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4717 float2367 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4718 float2368 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4719 LDBL[246] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=41d8   word=7   wl=18 address=0127
m4720 float2369 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4721 float2370 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4722 float2371 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4723 LDBL[55] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4724 LDBL[71] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4725 float2372 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4726 LDBL[103] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4727 LDBL[119] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4728 LDBL[135] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4729 float2373 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4730 float2374 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4731 float2375 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4732 float2376 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4733 float2377 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4734 LDBL[231] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4735 float2378 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a5e4   word=8   wl=18 address=0128
m4736 float2379 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4737 float2380 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4738 LDBL[40] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4739 float2381 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4740 float2382 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4741 LDBL[88] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4742 LDBL[104] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4743 LDBL[120] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4744 LDBL[136] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4745 float2383 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4746 LDBL[168] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4747 float2384 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4748 float2385 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4749 LDBL[216] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4750 float2386 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4751 LDBL[248] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f5b4   word=9   wl=18 address=0129
m4752 float2387 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4753 float2388 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4754 LDBL[41] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4755 float2389 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4756 LDBL[73] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4757 LDBL[89] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4758 float2390 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4759 LDBL[121] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4760 LDBL[137] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4761 float2391 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4762 LDBL[169] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4763 float2392 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4764 LDBL[201] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4765 LDBL[217] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4766 LDBL[233] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4767 LDBL[249] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0655   word=10   wl=18 address=012a
m4768 LDBL[10] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4769 float2393 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4770 LDBL[42] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4771 float2394 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4772 LDBL[74] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4773 float2395 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4774 LDBL[106] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4775 float2396 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4776 float2397 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4777 LDBL[154] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4778 LDBL[170] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4779 float2398 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4780 float2399 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4781 float2400 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4782 float2401 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4783 float2402 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=002f   word=11   wl=18 address=012b
m4784 LDBL[11] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4785 LDBL[27] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4786 LDBL[43] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4787 LDBL[59] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4788 float2403 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4789 LDBL[91] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4790 float2404 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4791 float2405 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4792 float2406 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4793 float2407 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4794 float2408 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4795 float2409 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4796 float2410 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4797 float2411 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4798 float2412 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4799 float2413 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6192   word=12   wl=18 address=012c
m4800 float2414 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4801 LDBL[28] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4802 float2415 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4803 float2416 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4804 LDBL[76] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4805 float2417 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4806 float2418 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4807 LDBL[124] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4808 LDBL[140] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4809 float2419 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4810 float2420 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4811 float2421 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4812 float2422 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4813 LDBL[220] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4814 LDBL[236] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4815 float2423 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d14d   word=13   wl=18 address=012d
m4816 LDBL[13] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4817 float2424 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4818 LDBL[45] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4819 LDBL[61] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4820 float2425 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4821 float2426 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4822 LDBL[109] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4823 float2427 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4824 LDBL[141] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4825 float2428 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4826 float2429 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4827 float2430 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4828 LDBL[205] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4829 float2431 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4830 LDBL[237] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4831 LDBL[253] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=831a   word=14   wl=18 address=012e
m4832 float2432 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4833 LDBL[30] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4834 float2433 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4835 LDBL[62] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4836 LDBL[78] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4837 float2434 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4838 float2435 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4839 float2436 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4840 LDBL[142] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4841 LDBL[158] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4842 float2437 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4843 float2438 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4844 float2439 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4845 float2440 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4846 float2441 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4847 LDBL[254] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fe36   word=15   wl=18 address=012f
m4848 float2442 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4849 LDBL[31] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4850 LDBL[47] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4851 float2443 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4852 LDBL[79] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4853 LDBL[95] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4854 float2444 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4855 float2445 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4856 float2446 LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4857 LDBL[159] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4858 LDBL[175] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4859 LDBL[191] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4860 LDBL[207] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4861 LDBL[223] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4862 LDBL[239] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4863 LDBL[255] LDWL[18] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4e04   word=0   wl=19 address=0130
m4864 float2447 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4865 float2448 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4866 LDBL[32] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4867 float2449 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4868 float2450 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4869 float2451 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4870 float2452 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4871 float2453 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4872 float2454 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4873 LDBL[144] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4874 LDBL[160] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4875 LDBL[176] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4876 float2455 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4877 float2456 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4878 LDBL[224] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4879 float2457 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b8e8   word=1   wl=19 address=0131
m4880 float2458 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4881 float2459 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4882 float2460 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4883 LDBL[49] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4884 float2461 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4885 LDBL[81] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4886 LDBL[97] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4887 LDBL[113] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4888 float2462 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4889 float2463 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4890 float2464 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4891 LDBL[177] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4892 LDBL[193] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4893 LDBL[209] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4894 float2465 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4895 LDBL[241] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f8a7   word=2   wl=19 address=0132
m4896 LDBL[2] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4897 LDBL[18] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4898 LDBL[34] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4899 float2466 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4900 float2467 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4901 LDBL[82] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4902 float2468 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4903 LDBL[114] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4904 float2469 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4905 float2470 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4906 float2471 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4907 LDBL[178] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4908 LDBL[194] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4909 LDBL[210] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4910 LDBL[226] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4911 LDBL[242] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9b16   word=3   wl=19 address=0133
m4912 float2472 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4913 LDBL[19] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4914 LDBL[35] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4915 float2473 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4916 LDBL[67] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4917 float2474 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4918 float2475 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4919 float2476 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4920 LDBL[131] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4921 LDBL[147] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4922 float2477 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4923 LDBL[179] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4924 LDBL[195] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4925 float2478 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4926 float2479 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4927 LDBL[243] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6384   word=4   wl=19 address=0134
m4928 float2480 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4929 float2481 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4930 LDBL[36] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4931 float2482 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4932 float2483 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4933 float2484 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4934 float2485 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4935 LDBL[116] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4936 LDBL[132] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4937 LDBL[148] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4938 float2486 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4939 float2487 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4940 float2488 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4941 LDBL[212] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4942 LDBL[228] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4943 float2489 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2590   word=5   wl=19 address=0135
m4944 float2490 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4945 float2491 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4946 float2492 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4947 float2493 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4948 LDBL[69] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4949 float2494 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4950 float2495 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4951 LDBL[117] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4952 LDBL[133] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4953 float2496 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4954 LDBL[165] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4955 float2497 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4956 float2498 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4957 LDBL[213] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4958 float2499 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4959 float2500 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0444   word=6   wl=19 address=0136
m4960 float2501 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4961 float2502 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4962 LDBL[38] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4963 float2503 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4964 float2504 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4965 float2505 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4966 LDBL[102] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4967 float2506 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4968 float2507 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4969 float2508 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4970 LDBL[166] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4971 float2509 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4972 float2510 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4973 float2511 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4974 float2512 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4975 float2513 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d380   word=7   wl=19 address=0137
m4976 float2514 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4977 float2515 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4978 float2516 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4979 float2517 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4980 float2518 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4981 float2519 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4982 float2520 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4983 LDBL[119] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4984 LDBL[135] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4985 LDBL[151] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4986 float2521 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4987 float2522 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4988 LDBL[199] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4989 float2523 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4990 LDBL[231] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4991 LDBL[247] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a81a   word=8   wl=19 address=0138
m4992 float2524 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4993 LDBL[24] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4994 float2525 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4995 LDBL[56] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4996 LDBL[72] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4997 float2526 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4998 float2527 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m4999 float2528 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5000 float2529 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5001 float2530 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5002 float2531 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5003 LDBL[184] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5004 float2532 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5005 LDBL[216] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5006 float2533 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5007 LDBL[248] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c924   word=9   wl=19 address=0139
m5008 float2534 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5009 float2535 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5010 LDBL[41] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5011 float2536 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5012 float2537 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5013 LDBL[89] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5014 float2538 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5015 float2539 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5016 LDBL[137] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5017 float2540 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5018 float2541 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5019 LDBL[185] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5020 float2542 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5021 float2543 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5022 LDBL[233] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5023 LDBL[249] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=868d   word=10   wl=19 address=013a
m5024 LDBL[10] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5025 float2544 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5026 LDBL[42] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5027 LDBL[58] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5028 float2545 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5029 float2546 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5030 float2547 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5031 LDBL[122] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5032 float2548 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5033 LDBL[154] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5034 LDBL[170] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5035 float2549 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5036 float2550 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5037 float2551 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5038 float2552 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5039 LDBL[250] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a086   word=11   wl=19 address=013b
m5040 float2553 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5041 LDBL[27] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5042 LDBL[43] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5043 float2554 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5044 float2555 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5045 float2556 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5046 float2557 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5047 LDBL[123] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5048 float2558 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5049 float2559 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5050 float2560 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5051 float2561 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5052 float2562 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5053 LDBL[219] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5054 float2563 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5055 LDBL[251] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a405   word=12   wl=19 address=013c
m5056 LDBL[12] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5057 float2564 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5058 LDBL[44] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5059 float2565 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5060 float2566 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5061 float2567 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5062 float2568 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5063 float2569 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5064 float2570 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5065 float2571 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5066 LDBL[172] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5067 float2572 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5068 float2573 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5069 LDBL[220] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5070 float2574 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5071 LDBL[252] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e37c   word=13   wl=19 address=013d
m5072 float2575 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5073 float2576 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5074 LDBL[45] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5075 LDBL[61] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5076 LDBL[77] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5077 LDBL[93] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5078 LDBL[109] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5079 float2577 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5080 LDBL[141] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5081 LDBL[157] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5082 float2578 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5083 float2579 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5084 float2580 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5085 LDBL[221] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5086 LDBL[237] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5087 LDBL[253] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=495f   word=14   wl=19 address=013e
m5088 LDBL[14] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5089 LDBL[30] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5090 LDBL[46] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5091 LDBL[62] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5092 LDBL[78] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5093 float2581 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5094 LDBL[110] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5095 float2582 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5096 LDBL[142] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5097 float2583 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5098 float2584 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5099 LDBL[190] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5100 float2585 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5101 float2586 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5102 LDBL[238] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5103 float2587 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=62ba   word=15   wl=19 address=013f
m5104 float2588 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5105 LDBL[31] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5106 float2589 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5107 LDBL[63] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5108 LDBL[79] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5109 LDBL[95] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5110 float2590 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5111 LDBL[127] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5112 float2591 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5113 LDBL[159] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5114 float2592 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5115 float2593 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5116 float2594 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5117 LDBL[223] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5118 LDBL[239] LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5119 float2595 LDWL[19] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ead5   word=0   wl=20 address=0140
m5120 LDBL[0] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5121 float2596 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5122 LDBL[32] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5123 float2597 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5124 LDBL[64] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5125 float2598 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5126 LDBL[96] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5127 LDBL[112] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5128 float2599 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5129 LDBL[144] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5130 float2600 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5131 LDBL[176] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5132 float2601 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5133 LDBL[208] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5134 LDBL[224] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5135 LDBL[240] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=443a   word=1   wl=20 address=0141
m5136 float2602 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5137 LDBL[17] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5138 float2603 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5139 LDBL[49] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5140 LDBL[65] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5141 LDBL[81] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5142 float2604 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5143 float2605 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5144 float2606 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5145 float2607 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5146 LDBL[161] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5147 float2608 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5148 float2609 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5149 float2610 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5150 LDBL[225] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5151 float2611 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7f45   word=2   wl=20 address=0142
m5152 LDBL[2] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5153 float2612 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5154 LDBL[34] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5155 float2613 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5156 float2614 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5157 float2615 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5158 LDBL[98] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5159 float2616 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5160 LDBL[130] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5161 LDBL[146] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5162 LDBL[162] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5163 LDBL[178] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5164 LDBL[194] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5165 LDBL[210] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5166 LDBL[226] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5167 float2617 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f437   word=3   wl=20 address=0143
m5168 LDBL[3] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5169 LDBL[19] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5170 LDBL[35] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5171 float2618 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5172 LDBL[67] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5173 LDBL[83] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5174 float2619 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5175 float2620 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5176 float2621 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5177 float2622 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5178 LDBL[163] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5179 float2623 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5180 LDBL[195] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5181 LDBL[211] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5182 LDBL[227] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5183 LDBL[243] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6b10   word=4   wl=20 address=0144
m5184 float2624 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5185 float2625 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5186 float2626 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5187 float2627 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5188 LDBL[68] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5189 float2628 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5190 float2629 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5191 float2630 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5192 LDBL[132] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5193 LDBL[148] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5194 float2631 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5195 LDBL[180] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5196 float2632 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5197 LDBL[212] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5198 LDBL[228] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5199 float2633 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=936a   word=5   wl=20 address=0145
m5200 float2634 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5201 LDBL[21] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5202 float2635 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5203 LDBL[53] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5204 float2636 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5205 LDBL[85] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5206 LDBL[101] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5207 float2637 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5208 LDBL[133] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5209 LDBL[149] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5210 float2638 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5211 float2639 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5212 LDBL[197] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5213 float2640 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5214 float2641 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5215 LDBL[245] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=073c   word=6   wl=20 address=0146
m5216 float2642 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5217 float2643 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5218 LDBL[38] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5219 LDBL[54] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5220 LDBL[70] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5221 LDBL[86] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5222 float2644 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5223 float2645 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5224 LDBL[134] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5225 LDBL[150] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5226 LDBL[166] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5227 float2646 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5228 float2647 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5229 float2648 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5230 float2649 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5231 float2650 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=679f   word=7   wl=20 address=0147
m5232 LDBL[7] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5233 LDBL[23] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5234 LDBL[39] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5235 LDBL[55] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5236 LDBL[71] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5237 float2651 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5238 float2652 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5239 LDBL[119] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5240 LDBL[135] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5241 LDBL[151] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5242 LDBL[167] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5243 float2653 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5244 float2654 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5245 LDBL[215] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5246 LDBL[231] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5247 float2655 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d96c   word=8   wl=20 address=0148
m5248 float2656 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5249 float2657 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5250 LDBL[40] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5251 LDBL[56] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5252 float2658 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5253 LDBL[88] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5254 LDBL[104] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5255 float2659 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5256 LDBL[136] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5257 float2660 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5258 float2661 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5259 LDBL[184] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5260 LDBL[200] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5261 float2662 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5262 LDBL[232] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5263 LDBL[248] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9cf8   word=9   wl=20 address=0149
m5264 float2663 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5265 float2664 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5266 float2665 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5267 LDBL[57] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5268 LDBL[73] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5269 LDBL[89] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5270 LDBL[105] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5271 LDBL[121] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5272 float2666 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5273 float2667 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5274 LDBL[169] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5275 LDBL[185] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5276 LDBL[201] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5277 float2668 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5278 float2669 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5279 LDBL[249] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a298   word=10   wl=20 address=014a
m5280 float2670 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5281 float2671 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5282 float2672 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5283 LDBL[58] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5284 LDBL[74] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5285 float2673 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5286 float2674 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5287 LDBL[122] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5288 float2675 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5289 LDBL[154] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5290 float2676 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5291 float2677 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5292 float2678 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5293 LDBL[218] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5294 float2679 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5295 LDBL[250] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=dab8   word=11   wl=20 address=014b
m5296 float2680 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5297 float2681 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5298 float2682 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5299 LDBL[59] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5300 LDBL[75] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5301 LDBL[91] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5302 float2683 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5303 LDBL[123] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5304 float2684 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5305 LDBL[155] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5306 float2685 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5307 LDBL[187] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5308 LDBL[203] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5309 float2686 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5310 LDBL[235] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5311 LDBL[251] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=bd46   word=12   wl=20 address=014c
m5312 float2687 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5313 LDBL[28] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5314 LDBL[44] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5315 float2688 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5316 float2689 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5317 float2690 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5318 LDBL[108] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5319 float2691 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5320 LDBL[140] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5321 float2692 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5322 LDBL[172] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5323 LDBL[188] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5324 LDBL[204] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5325 LDBL[220] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5326 float2693 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5327 LDBL[252] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2581   word=13   wl=20 address=014d
m5328 LDBL[13] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5329 float2694 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5330 float2695 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5331 float2696 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5332 float2697 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5333 float2698 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5334 float2699 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5335 LDBL[125] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5336 LDBL[141] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5337 float2700 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5338 LDBL[173] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5339 float2701 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5340 float2702 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5341 LDBL[221] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5342 float2703 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5343 float2704 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=659c   word=14   wl=20 address=014e
m5344 float2705 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5345 float2706 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5346 LDBL[46] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5347 LDBL[62] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5348 LDBL[78] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5349 float2707 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5350 float2708 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5351 LDBL[126] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5352 LDBL[142] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5353 float2709 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5354 LDBL[174] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5355 float2710 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5356 float2711 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5357 LDBL[222] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5358 LDBL[238] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5359 float2712 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ee41   word=15   wl=20 address=014f
m5360 LDBL[15] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5361 float2713 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5362 float2714 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5363 float2715 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5364 float2716 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5365 float2717 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5366 LDBL[111] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5367 float2718 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5368 float2719 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5369 LDBL[159] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5370 LDBL[175] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5371 LDBL[191] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5372 float2720 LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5373 LDBL[223] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5374 LDBL[239] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5375 LDBL[255] LDWL[20] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4b15   word=0   wl=21 address=0150
m5376 LDBL[0] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5377 float2721 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5378 LDBL[32] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5379 float2722 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5380 LDBL[64] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5381 float2723 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5382 float2724 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5383 float2725 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5384 LDBL[128] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5385 LDBL[144] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5386 float2726 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5387 LDBL[176] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5388 float2727 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5389 float2728 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5390 LDBL[224] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5391 float2729 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=cdb3   word=1   wl=21 address=0151
m5392 LDBL[1] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5393 LDBL[17] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5394 float2730 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5395 float2731 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5396 LDBL[65] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5397 LDBL[81] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5398 float2732 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5399 LDBL[113] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5400 LDBL[129] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5401 float2733 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5402 LDBL[161] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5403 LDBL[177] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5404 float2734 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5405 float2735 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5406 LDBL[225] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5407 LDBL[241] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=882f   word=2   wl=21 address=0152
m5408 LDBL[2] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5409 LDBL[18] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5410 LDBL[34] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5411 LDBL[50] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5412 float2736 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5413 LDBL[82] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5414 float2737 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5415 float2738 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5416 float2739 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5417 float2740 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5418 float2741 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5419 LDBL[178] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5420 float2742 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5421 float2743 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5422 float2744 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5423 LDBL[242] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=867f   word=3   wl=21 address=0153
m5424 LDBL[3] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5425 LDBL[19] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5426 LDBL[35] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5427 LDBL[51] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5428 LDBL[67] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5429 LDBL[83] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5430 LDBL[99] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5431 float2745 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5432 float2746 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5433 LDBL[147] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5434 LDBL[163] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5435 float2747 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5436 float2748 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5437 float2749 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5438 float2750 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5439 LDBL[243] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=275d   word=4   wl=21 address=0154
m5440 LDBL[4] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5441 float2751 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5442 LDBL[36] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5443 LDBL[52] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5444 LDBL[68] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5445 float2752 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5446 LDBL[100] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5447 float2753 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5448 LDBL[132] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5449 LDBL[148] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5450 LDBL[164] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5451 float2754 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5452 float2755 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5453 LDBL[212] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5454 float2756 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5455 float2757 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6750   word=5   wl=21 address=0155
m5456 float2758 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5457 float2759 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5458 float2760 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5459 float2761 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5460 LDBL[69] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5461 float2762 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5462 LDBL[101] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5463 float2763 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5464 LDBL[133] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5465 LDBL[149] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5466 LDBL[165] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5467 float2764 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5468 float2765 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5469 LDBL[213] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5470 LDBL[229] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5471 float2766 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=16d1   word=6   wl=21 address=0156
m5472 LDBL[6] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5473 float2767 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5474 float2768 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5475 float2769 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5476 LDBL[70] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5477 float2770 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5478 LDBL[102] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5479 LDBL[118] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5480 float2771 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5481 LDBL[150] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5482 LDBL[166] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5483 float2772 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5484 LDBL[198] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5485 float2773 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5486 float2774 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5487 float2775 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1adb   word=7   wl=21 address=0157
m5488 LDBL[7] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5489 LDBL[23] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5490 float2776 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5491 LDBL[55] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5492 LDBL[71] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5493 float2777 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5494 LDBL[103] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5495 LDBL[119] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5496 float2778 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5497 LDBL[151] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5498 float2779 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5499 LDBL[183] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5500 LDBL[199] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5501 float2780 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5502 float2781 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5503 float2782 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2551   word=8   wl=21 address=0158
m5504 LDBL[8] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5505 float2783 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5506 float2784 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5507 float2785 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5508 LDBL[72] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5509 float2786 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5510 LDBL[104] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5511 float2787 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5512 LDBL[136] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5513 float2788 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5514 LDBL[168] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5515 float2789 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5516 float2790 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5517 LDBL[216] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5518 float2791 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5519 float2792 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=cf78   word=9   wl=21 address=0159
m5520 float2793 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5521 float2794 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5522 float2795 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5523 LDBL[57] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5524 LDBL[73] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5525 LDBL[89] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5526 LDBL[105] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5527 float2796 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5528 LDBL[137] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5529 LDBL[153] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5530 LDBL[169] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5531 LDBL[185] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5532 float2797 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5533 float2798 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5534 LDBL[233] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5535 LDBL[249] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a8ed   word=10   wl=21 address=015a
m5536 LDBL[10] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5537 float2799 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5538 LDBL[42] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5539 LDBL[58] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5540 float2800 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5541 LDBL[90] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5542 LDBL[106] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5543 LDBL[122] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5544 float2801 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5545 float2802 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5546 float2803 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5547 LDBL[186] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5548 float2804 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5549 LDBL[218] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5550 float2805 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5551 LDBL[250] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f24f   word=11   wl=21 address=015b
m5552 LDBL[11] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5553 LDBL[27] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5554 LDBL[43] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5555 LDBL[59] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5556 float2806 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5557 float2807 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5558 LDBL[107] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5559 float2808 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5560 float2809 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5561 LDBL[155] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5562 float2810 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5563 float2811 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5564 LDBL[203] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5565 LDBL[219] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5566 LDBL[235] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5567 LDBL[251] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fb0b   word=12   wl=21 address=015c
m5568 LDBL[12] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5569 LDBL[28] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5570 float2812 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5571 LDBL[60] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5572 float2813 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5573 float2814 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5574 float2815 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5575 float2816 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5576 LDBL[140] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5577 LDBL[156] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5578 float2817 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5579 LDBL[188] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5580 LDBL[204] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5581 LDBL[220] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5582 LDBL[236] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5583 LDBL[252] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1af8   word=13   wl=21 address=015d
m5584 float2818 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5585 float2819 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5586 float2820 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5587 LDBL[61] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5588 LDBL[77] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5589 LDBL[93] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5590 LDBL[109] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5591 LDBL[125] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5592 float2821 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5593 LDBL[157] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5594 float2822 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5595 LDBL[189] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5596 LDBL[205] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5597 float2823 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5598 float2824 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5599 float2825 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=193b   word=14   wl=21 address=015e
m5600 LDBL[14] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5601 LDBL[30] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5602 float2826 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5603 LDBL[62] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5604 LDBL[78] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5605 LDBL[94] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5606 float2827 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5607 float2828 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5608 LDBL[142] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5609 float2829 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5610 float2830 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5611 LDBL[190] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5612 LDBL[206] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5613 float2831 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5614 float2832 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5615 float2833 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c671   word=15   wl=21 address=015f
m5616 LDBL[15] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5617 float2834 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5618 float2835 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5619 float2836 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5620 LDBL[79] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5621 LDBL[95] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5622 LDBL[111] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5623 float2837 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5624 float2838 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5625 LDBL[159] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5626 LDBL[175] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5627 float2839 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5628 float2840 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5629 float2841 LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5630 LDBL[239] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5631 LDBL[255] LDWL[21] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4b8c   word=0   wl=22 address=0160
m5632 float2842 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5633 float2843 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5634 LDBL[32] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5635 LDBL[48] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5636 float2844 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5637 float2845 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5638 float2846 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5639 LDBL[112] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5640 LDBL[128] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5641 LDBL[144] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5642 float2847 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5643 LDBL[176] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5644 float2848 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5645 float2849 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5646 LDBL[224] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5647 float2850 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1af9   word=1   wl=22 address=0161
m5648 LDBL[1] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5649 float2851 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5650 float2852 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5651 LDBL[49] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5652 LDBL[65] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5653 LDBL[81] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5654 LDBL[97] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5655 LDBL[113] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5656 float2853 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5657 LDBL[145] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5658 float2854 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5659 LDBL[177] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5660 LDBL[193] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5661 float2855 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5662 float2856 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5663 float2857 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ad25   word=2   wl=22 address=0162
m5664 LDBL[2] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5665 float2858 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5666 LDBL[34] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5667 float2859 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5668 float2860 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5669 LDBL[82] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5670 float2861 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5671 float2862 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5672 LDBL[130] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5673 float2863 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5674 LDBL[162] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5675 LDBL[178] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5676 float2864 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5677 LDBL[210] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5678 float2865 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5679 LDBL[242] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7709   word=3   wl=22 address=0163
m5680 LDBL[3] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5681 float2866 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5682 float2867 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5683 LDBL[51] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5684 float2868 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5685 float2869 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5686 float2870 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5687 float2871 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5688 LDBL[131] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5689 LDBL[147] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5690 LDBL[163] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5691 float2872 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5692 LDBL[195] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5693 LDBL[211] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5694 LDBL[227] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5695 float2873 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a3f9   word=4   wl=22 address=0164
m5696 LDBL[4] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5697 float2874 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5698 float2875 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5699 LDBL[52] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5700 LDBL[68] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5701 LDBL[84] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5702 LDBL[100] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5703 LDBL[116] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5704 LDBL[132] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5705 LDBL[148] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5706 float2876 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5707 float2877 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5708 float2878 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5709 LDBL[212] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5710 float2879 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5711 LDBL[244] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=43c6   word=5   wl=22 address=0165
m5712 float2880 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5713 LDBL[21] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5714 LDBL[37] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5715 float2881 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5716 float2882 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5717 float2883 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5718 LDBL[101] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5719 LDBL[117] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5720 LDBL[133] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5721 LDBL[149] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5722 float2884 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5723 float2885 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5724 float2886 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5725 float2887 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5726 LDBL[229] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5727 float2888 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=767a   word=6   wl=22 address=0166
m5728 float2889 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5729 LDBL[22] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5730 float2890 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5731 LDBL[54] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5732 LDBL[70] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5733 LDBL[86] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5734 LDBL[102] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5735 float2891 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5736 float2892 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5737 LDBL[150] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5738 LDBL[166] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5739 float2893 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5740 LDBL[198] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5741 LDBL[214] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5742 LDBL[230] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5743 float2894 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=36f0   word=7   wl=22 address=0167
m5744 float2895 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5745 float2896 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5746 float2897 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5747 float2898 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5748 LDBL[71] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5749 LDBL[87] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5750 LDBL[103] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5751 LDBL[119] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5752 float2899 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5753 LDBL[151] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5754 LDBL[167] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5755 float2900 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5756 LDBL[199] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5757 LDBL[215] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5758 float2901 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5759 float2902 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e07f   word=8   wl=22 address=0168
m5760 LDBL[8] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5761 LDBL[24] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5762 LDBL[40] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5763 LDBL[56] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5764 LDBL[72] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5765 LDBL[88] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5766 LDBL[104] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5767 float2903 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5768 float2904 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5769 float2905 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5770 float2906 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5771 float2907 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5772 float2908 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5773 LDBL[216] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5774 LDBL[232] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5775 LDBL[248] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1e5f   word=9   wl=22 address=0169
m5776 LDBL[9] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5777 LDBL[25] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5778 LDBL[41] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5779 LDBL[57] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5780 LDBL[73] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5781 float2909 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5782 LDBL[105] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5783 float2910 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5784 float2911 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5785 LDBL[153] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5786 LDBL[169] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5787 LDBL[185] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5788 LDBL[201] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5789 float2912 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5790 float2913 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5791 float2914 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=317c   word=10   wl=22 address=016a
m5792 float2915 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5793 float2916 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5794 LDBL[42] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5795 LDBL[58] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5796 LDBL[74] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5797 LDBL[90] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5798 LDBL[106] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5799 float2917 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5800 LDBL[138] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5801 float2918 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5802 float2919 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5803 float2920 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5804 LDBL[202] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5805 LDBL[218] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5806 float2921 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5807 float2922 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3356   word=11   wl=22 address=016b
m5808 float2923 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5809 LDBL[27] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5810 LDBL[43] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5811 float2924 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5812 LDBL[75] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5813 float2925 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5814 LDBL[107] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5815 float2926 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5816 LDBL[139] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5817 LDBL[155] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5818 float2927 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5819 float2928 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5820 LDBL[203] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5821 LDBL[219] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5822 float2929 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5823 float2930 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f2b5   word=12   wl=22 address=016c
m5824 LDBL[12] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5825 float2931 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5826 LDBL[44] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5827 float2932 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5828 LDBL[76] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5829 LDBL[92] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5830 float2933 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5831 LDBL[124] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5832 float2934 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5833 LDBL[156] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5834 float2935 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5835 float2936 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5836 LDBL[204] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5837 LDBL[220] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5838 LDBL[236] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5839 LDBL[252] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5dc0   word=13   wl=22 address=016d
m5840 float2937 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5841 float2938 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5842 float2939 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5843 float2940 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5844 float2941 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5845 float2942 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5846 LDBL[109] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5847 LDBL[125] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5848 LDBL[141] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5849 float2943 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5850 LDBL[173] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5851 LDBL[189] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5852 LDBL[205] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5853 float2944 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5854 LDBL[237] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5855 float2945 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5193   word=14   wl=22 address=016e
m5856 LDBL[14] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5857 LDBL[30] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5858 float2946 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5859 float2947 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5860 LDBL[78] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5861 float2948 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5862 float2949 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5863 LDBL[126] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5864 LDBL[142] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5865 float2950 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5866 float2951 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5867 float2952 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5868 LDBL[206] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5869 float2953 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5870 LDBL[238] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5871 float2954 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5e9f   word=15   wl=22 address=016f
m5872 LDBL[15] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5873 LDBL[31] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5874 LDBL[47] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5875 LDBL[63] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5876 LDBL[79] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5877 float2955 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5878 float2956 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5879 LDBL[127] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5880 float2957 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5881 LDBL[159] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5882 LDBL[175] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5883 LDBL[191] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5884 LDBL[207] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5885 float2958 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5886 LDBL[239] LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5887 float2959 LDWL[22] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8b4e   word=0   wl=23 address=0170
m5888 float2960 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5889 LDBL[16] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5890 LDBL[32] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5891 LDBL[48] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5892 float2961 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5893 float2962 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5894 LDBL[96] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5895 float2963 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5896 LDBL[128] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5897 LDBL[144] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5898 float2964 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5899 LDBL[176] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5900 float2965 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5901 float2966 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5902 float2967 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5903 LDBL[240] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1c79   word=1   wl=23 address=0171
m5904 LDBL[1] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5905 float2968 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5906 float2969 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5907 LDBL[49] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5908 LDBL[65] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5909 LDBL[81] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5910 LDBL[97] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5911 float2970 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5912 float2971 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5913 float2972 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5914 LDBL[161] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5915 LDBL[177] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5916 LDBL[193] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5917 float2973 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5918 float2974 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5919 float2975 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e63c   word=2   wl=23 address=0172
m5920 float2976 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5921 float2977 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5922 LDBL[34] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5923 LDBL[50] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5924 LDBL[66] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5925 LDBL[82] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5926 float2978 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5927 float2979 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5928 float2980 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5929 LDBL[146] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5930 LDBL[162] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5931 float2981 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5932 float2982 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5933 LDBL[210] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5934 LDBL[226] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5935 LDBL[242] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5899   word=3   wl=23 address=0173
m5936 LDBL[3] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5937 float2983 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5938 float2984 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5939 LDBL[51] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5940 LDBL[67] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5941 float2985 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5942 float2986 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5943 LDBL[115] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5944 float2987 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5945 float2988 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5946 float2989 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5947 LDBL[179] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5948 LDBL[195] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5949 float2990 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5950 LDBL[227] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5951 float2991 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5f20   word=4   wl=23 address=0174
m5952 float2992 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5953 float2993 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5954 float2994 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5955 float2995 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5956 float2996 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5957 LDBL[84] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5958 float2997 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5959 float2998 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5960 LDBL[132] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5961 LDBL[148] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5962 LDBL[164] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5963 LDBL[180] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5964 LDBL[196] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5965 float2999 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5966 LDBL[228] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5967 float3000 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a5a8   word=5   wl=23 address=0175
m5968 float3001 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5969 float3002 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5970 float3003 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5971 LDBL[53] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5972 float3004 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5973 LDBL[85] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5974 float3005 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5975 LDBL[117] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5976 LDBL[133] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5977 float3006 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5978 LDBL[165] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5979 float3007 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5980 float3008 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5981 LDBL[213] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5982 float3009 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5983 LDBL[245] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8391   word=6   wl=23 address=0176
m5984 LDBL[6] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5985 float3010 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5986 float3011 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5987 float3012 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5988 LDBL[70] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5989 float3013 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5990 float3014 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5991 LDBL[118] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5992 LDBL[134] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5993 LDBL[150] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5994 float3015 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5995 float3016 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5996 float3017 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5997 float3018 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5998 float3019 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m5999 LDBL[246] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=94a9   word=7   wl=23 address=0177
m6000 LDBL[7] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6001 float3020 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6002 float3021 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6003 LDBL[55] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6004 float3022 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6005 LDBL[87] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6006 float3023 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6007 LDBL[119] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6008 float3024 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6009 float3025 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6010 LDBL[167] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6011 float3026 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6012 LDBL[199] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6013 float3027 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6014 float3028 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6015 LDBL[247] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5dd9   word=8   wl=23 address=0178
m6016 LDBL[8] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6017 float3029 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6018 float3030 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6019 LDBL[56] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6020 LDBL[72] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6021 float3031 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6022 LDBL[104] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6023 LDBL[120] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6024 LDBL[136] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6025 float3032 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6026 LDBL[168] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6027 LDBL[184] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6028 LDBL[200] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6029 float3033 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6030 LDBL[232] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6031 float3034 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d60a   word=9   wl=23 address=0179
m6032 float3035 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6033 LDBL[25] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6034 float3036 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6035 LDBL[57] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6036 float3037 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6037 float3038 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6038 float3039 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6039 float3040 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6040 float3041 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6041 LDBL[153] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6042 LDBL[169] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6043 float3042 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6044 LDBL[201] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6045 float3043 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6046 LDBL[233] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6047 LDBL[249] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b4b9   word=10   wl=23 address=017a
m6048 LDBL[10] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6049 float3044 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6050 float3045 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6051 LDBL[58] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6052 LDBL[74] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6053 LDBL[90] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6054 float3046 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6055 LDBL[122] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6056 float3047 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6057 float3048 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6058 LDBL[170] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6059 float3049 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6060 LDBL[202] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6061 LDBL[218] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6062 float3050 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6063 LDBL[250] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=65f1   word=11   wl=23 address=017b
m6064 LDBL[11] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6065 float3051 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6066 float3052 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6067 float3053 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6068 LDBL[75] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6069 LDBL[91] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6070 LDBL[107] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6071 LDBL[123] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6072 LDBL[139] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6073 float3054 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6074 LDBL[171] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6075 float3055 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6076 float3056 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6077 LDBL[219] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6078 LDBL[235] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6079 float3057 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b2fd   word=12   wl=23 address=017c
m6080 LDBL[12] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6081 float3058 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6082 LDBL[44] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6083 LDBL[60] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6084 LDBL[76] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6085 LDBL[92] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6086 LDBL[108] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6087 LDBL[124] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6088 float3059 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6089 LDBL[156] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6090 float3060 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6091 float3061 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6092 LDBL[204] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6093 LDBL[220] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6094 float3062 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6095 LDBL[252] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2111   word=13   wl=23 address=017d
m6096 LDBL[13] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6097 float3063 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6098 float3064 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6099 float3065 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6100 LDBL[77] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6101 float3066 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6102 float3067 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6103 float3068 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6104 LDBL[141] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6105 float3069 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6106 float3070 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6107 float3071 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6108 float3072 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6109 LDBL[221] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6110 float3073 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6111 float3074 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2dd6   word=14   wl=23 address=017e
m6112 float3075 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6113 LDBL[30] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6114 LDBL[46] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6115 float3076 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6116 LDBL[78] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6117 float3077 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6118 LDBL[110] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6119 LDBL[126] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6120 LDBL[142] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6121 float3078 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6122 LDBL[174] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6123 LDBL[190] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6124 float3079 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6125 LDBL[222] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6126 float3080 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6127 float3081 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=620f   word=15   wl=23 address=017f
m6128 LDBL[15] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6129 LDBL[31] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6130 LDBL[47] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6131 LDBL[63] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6132 float3082 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6133 float3083 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6134 float3084 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6135 float3085 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6136 float3086 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6137 LDBL[159] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6138 float3087 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6139 float3088 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6140 float3089 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6141 LDBL[223] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6142 LDBL[239] LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6143 float3090 LDWL[23] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5bb5   word=0   wl=24 address=0180
m6144 LDBL[0] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6145 float3091 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6146 LDBL[32] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6147 float3092 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6148 LDBL[64] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6149 LDBL[80] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6150 float3093 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6151 LDBL[112] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6152 LDBL[128] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6153 LDBL[144] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6154 float3094 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6155 LDBL[176] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6156 LDBL[192] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6157 float3095 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6158 LDBL[224] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6159 float3096 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3c53   word=1   wl=24 address=0181
m6160 LDBL[1] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6161 LDBL[17] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6162 float3097 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6163 float3098 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6164 LDBL[65] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6165 float3099 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6166 LDBL[97] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6167 float3100 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6168 float3101 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6169 float3102 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6170 LDBL[161] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6171 LDBL[177] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6172 LDBL[193] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6173 LDBL[209] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6174 float3103 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6175 float3104 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9bf7   word=2   wl=24 address=0182
m6176 LDBL[2] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6177 LDBL[18] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6178 LDBL[34] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6179 float3105 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6180 LDBL[66] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6181 LDBL[82] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6182 LDBL[98] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6183 LDBL[114] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6184 LDBL[130] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6185 LDBL[146] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6186 float3106 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6187 LDBL[178] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6188 LDBL[194] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6189 float3107 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6190 float3108 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6191 LDBL[242] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fb13   word=3   wl=24 address=0183
m6192 LDBL[3] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6193 LDBL[19] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6194 float3109 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6195 float3110 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6196 LDBL[67] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6197 float3111 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6198 float3112 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6199 float3113 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6200 LDBL[131] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6201 LDBL[147] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6202 float3114 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6203 LDBL[179] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6204 LDBL[195] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6205 LDBL[211] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6206 LDBL[227] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6207 LDBL[243] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6cde   word=4   wl=24 address=0184
m6208 float3115 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6209 LDBL[20] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6210 LDBL[36] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6211 LDBL[52] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6212 LDBL[68] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6213 float3116 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6214 LDBL[100] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6215 LDBL[116] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6216 float3117 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6217 float3118 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6218 LDBL[164] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6219 LDBL[180] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6220 float3119 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6221 LDBL[212] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6222 LDBL[228] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6223 float3120 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=448c   word=5   wl=24 address=0185
m6224 float3121 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6225 float3122 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6226 LDBL[37] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6227 LDBL[53] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6228 float3123 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6229 float3124 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6230 float3125 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6231 LDBL[117] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6232 float3126 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6233 float3127 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6234 LDBL[165] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6235 float3128 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6236 float3129 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6237 float3130 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6238 LDBL[229] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6239 float3131 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ebbd   word=6   wl=24 address=0186
m6240 LDBL[6] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6241 float3132 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6242 LDBL[38] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6243 LDBL[54] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6244 LDBL[70] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6245 LDBL[86] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6246 float3133 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6247 LDBL[118] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6248 LDBL[134] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6249 LDBL[150] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6250 float3134 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6251 LDBL[182] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6252 float3135 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6253 LDBL[214] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6254 LDBL[230] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6255 LDBL[246] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=193a   word=7   wl=24 address=0187
m6256 float3136 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6257 LDBL[23] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6258 float3137 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6259 LDBL[55] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6260 LDBL[71] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6261 LDBL[87] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6262 float3138 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6263 float3139 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6264 LDBL[135] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6265 float3140 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6266 float3141 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6267 LDBL[183] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6268 LDBL[199] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6269 float3142 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6270 float3143 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6271 float3144 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=79f7   word=8   wl=24 address=0188
m6272 LDBL[8] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6273 LDBL[24] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6274 LDBL[40] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6275 float3145 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6276 LDBL[72] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6277 LDBL[88] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6278 LDBL[104] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6279 LDBL[120] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6280 LDBL[136] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6281 float3146 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6282 float3147 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6283 LDBL[184] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6284 LDBL[200] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6285 LDBL[216] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6286 LDBL[232] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6287 float3148 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8c3b   word=9   wl=24 address=0189
m6288 LDBL[9] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6289 LDBL[25] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6290 float3149 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6291 LDBL[57] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6292 LDBL[73] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6293 LDBL[89] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6294 float3150 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6295 float3151 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6296 float3152 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6297 float3153 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6298 LDBL[169] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6299 LDBL[185] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6300 float3154 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6301 float3155 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6302 float3156 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6303 LDBL[249] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a46e   word=10   wl=24 address=018a
m6304 float3157 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6305 LDBL[26] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6306 LDBL[42] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6307 LDBL[58] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6308 float3158 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6309 LDBL[90] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6310 LDBL[106] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6311 float3159 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6312 float3160 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6313 float3161 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6314 LDBL[170] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6315 float3162 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6316 float3163 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6317 LDBL[218] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6318 float3164 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6319 LDBL[250] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4cbd   word=11   wl=24 address=018b
m6320 LDBL[11] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6321 float3165 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6322 LDBL[43] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6323 LDBL[59] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6324 LDBL[75] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6325 LDBL[91] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6326 float3166 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6327 LDBL[123] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6328 float3167 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6329 float3168 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6330 LDBL[171] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6331 LDBL[187] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6332 float3169 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6333 float3170 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6334 LDBL[235] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6335 float3171 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9bb3   word=12   wl=24 address=018c
m6336 LDBL[12] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6337 LDBL[28] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6338 float3172 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6339 float3173 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6340 LDBL[76] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6341 LDBL[92] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6342 float3174 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6343 LDBL[124] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6344 LDBL[140] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6345 LDBL[156] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6346 float3175 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6347 LDBL[188] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6348 LDBL[204] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6349 float3176 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6350 float3177 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6351 LDBL[252] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4618   word=13   wl=24 address=018d
m6352 float3178 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6353 float3179 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6354 float3180 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6355 LDBL[61] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6356 LDBL[77] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6357 float3181 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6358 float3182 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6359 float3183 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6360 float3184 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6361 LDBL[157] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6362 LDBL[173] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6363 float3185 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6364 float3186 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6365 float3187 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6366 LDBL[237] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6367 float3188 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6a9e   word=14   wl=24 address=018e
m6368 float3189 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6369 LDBL[30] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6370 LDBL[46] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6371 LDBL[62] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6372 LDBL[78] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6373 float3190 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6374 float3191 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6375 LDBL[126] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6376 float3192 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6377 LDBL[158] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6378 float3193 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6379 LDBL[190] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6380 float3194 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6381 LDBL[222] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6382 LDBL[238] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6383 float3195 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3ae1   word=15   wl=24 address=018f
m6384 LDBL[15] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6385 float3196 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6386 float3197 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6387 float3198 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6388 float3199 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6389 LDBL[95] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6390 LDBL[111] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6391 LDBL[127] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6392 float3200 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6393 LDBL[159] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6394 float3201 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6395 LDBL[191] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6396 LDBL[207] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6397 LDBL[223] LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6398 float3202 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6399 float3203 LDWL[24] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=857b   word=0   wl=25 address=0190
m6400 LDBL[0] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6401 LDBL[16] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6402 float3204 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6403 LDBL[48] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6404 LDBL[64] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6405 LDBL[80] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6406 LDBL[96] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6407 float3205 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6408 LDBL[128] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6409 float3206 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6410 LDBL[160] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6411 float3207 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6412 float3208 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6413 float3209 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6414 float3210 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6415 LDBL[240] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b916   word=1   wl=25 address=0191
m6416 float3211 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6417 LDBL[17] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6418 LDBL[33] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6419 float3212 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6420 LDBL[65] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6421 float3213 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6422 float3214 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6423 float3215 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6424 LDBL[129] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6425 float3216 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6426 float3217 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6427 LDBL[177] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6428 LDBL[193] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6429 LDBL[209] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6430 float3218 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6431 LDBL[241] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c27d   word=2   wl=25 address=0192
m6432 LDBL[2] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6433 float3219 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6434 LDBL[34] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6435 LDBL[50] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6436 LDBL[66] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6437 LDBL[82] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6438 LDBL[98] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6439 float3220 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6440 float3221 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6441 LDBL[146] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6442 float3222 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6443 float3223 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6444 float3224 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6445 float3225 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6446 LDBL[226] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6447 LDBL[242] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d077   word=3   wl=25 address=0193
m6448 LDBL[3] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6449 LDBL[19] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6450 LDBL[35] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6451 float3226 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6452 LDBL[67] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6453 LDBL[83] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6454 LDBL[99] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6455 float3227 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6456 float3228 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6457 float3229 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6458 float3230 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6459 float3231 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6460 LDBL[195] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6461 float3232 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6462 LDBL[227] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6463 LDBL[243] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=74e9   word=4   wl=25 address=0194
m6464 LDBL[4] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6465 float3233 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6466 float3234 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6467 LDBL[52] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6468 float3235 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6469 LDBL[84] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6470 LDBL[100] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6471 LDBL[116] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6472 float3236 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6473 float3237 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6474 LDBL[164] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6475 float3238 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6476 LDBL[196] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6477 LDBL[212] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6478 LDBL[228] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6479 float3239 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7ced   word=5   wl=25 address=0195
m6480 LDBL[5] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6481 float3240 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6482 LDBL[37] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6483 LDBL[53] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6484 float3241 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6485 LDBL[85] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6486 LDBL[101] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6487 LDBL[117] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6488 float3242 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6489 float3243 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6490 LDBL[165] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6491 LDBL[181] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6492 LDBL[197] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6493 LDBL[213] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6494 LDBL[229] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6495 float3244 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=dd9c   word=6   wl=25 address=0196
m6496 float3245 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6497 float3246 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6498 LDBL[38] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6499 LDBL[54] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6500 LDBL[70] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6501 float3247 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6502 float3248 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6503 LDBL[118] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6504 LDBL[134] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6505 float3249 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6506 LDBL[166] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6507 LDBL[182] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6508 LDBL[198] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6509 float3250 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6510 LDBL[230] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6511 LDBL[246] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b78a   word=7   wl=25 address=0197
m6512 float3251 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6513 LDBL[23] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6514 float3252 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6515 LDBL[55] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6516 float3253 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6517 float3254 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6518 float3255 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6519 LDBL[119] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6520 LDBL[135] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6521 LDBL[151] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6522 LDBL[167] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6523 float3256 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6524 LDBL[199] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6525 LDBL[215] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6526 float3257 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6527 LDBL[247] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=20b6   word=8   wl=25 address=0198
m6528 float3258 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6529 LDBL[24] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6530 LDBL[40] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6531 float3259 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6532 LDBL[72] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6533 LDBL[88] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6534 float3260 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6535 LDBL[120] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6536 float3261 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6537 float3262 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6538 float3263 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6539 float3264 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6540 float3265 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6541 LDBL[216] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6542 float3266 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6543 float3267 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1c0f   word=9   wl=25 address=0199
m6544 LDBL[9] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6545 LDBL[25] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6546 LDBL[41] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6547 LDBL[57] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6548 float3268 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6549 float3269 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6550 float3270 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6551 float3271 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6552 float3272 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6553 float3273 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6554 LDBL[169] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6555 LDBL[185] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6556 LDBL[201] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6557 float3274 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6558 float3275 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6559 float3276 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=43d6   word=10   wl=25 address=019a
m6560 float3277 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6561 LDBL[26] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6562 LDBL[42] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6563 float3278 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6564 LDBL[74] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6565 float3279 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6566 LDBL[106] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6567 LDBL[122] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6568 LDBL[138] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6569 LDBL[154] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6570 float3280 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6571 float3281 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6572 float3282 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6573 float3283 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6574 LDBL[234] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6575 float3284 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1ae5   word=11   wl=25 address=019b
m6576 LDBL[11] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6577 float3285 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6578 LDBL[43] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6579 float3286 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6580 float3287 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6581 LDBL[91] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6582 LDBL[107] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6583 LDBL[123] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6584 float3288 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6585 LDBL[155] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6586 float3289 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6587 LDBL[187] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6588 LDBL[203] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6589 float3290 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6590 float3291 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6591 float3292 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8fab   word=12   wl=25 address=019c
m6592 LDBL[12] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6593 LDBL[28] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6594 float3293 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6595 LDBL[60] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6596 float3294 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6597 LDBL[92] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6598 float3295 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6599 LDBL[124] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6600 LDBL[140] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6601 LDBL[156] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6602 LDBL[172] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6603 LDBL[188] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6604 float3296 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6605 float3297 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6606 float3298 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6607 LDBL[252] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3d72   word=13   wl=25 address=019d
m6608 float3299 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6609 LDBL[29] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6610 float3300 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6611 float3301 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6612 LDBL[77] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6613 LDBL[93] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6614 LDBL[109] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6615 float3302 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6616 LDBL[141] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6617 float3303 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6618 LDBL[173] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6619 LDBL[189] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6620 LDBL[205] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6621 LDBL[221] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6622 float3304 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6623 float3305 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=05a0   word=14   wl=25 address=019e
m6624 float3306 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6625 float3307 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6626 float3308 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6627 float3309 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6628 float3310 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6629 LDBL[94] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6630 float3311 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6631 LDBL[126] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6632 LDBL[142] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6633 float3312 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6634 LDBL[174] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6635 float3313 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6636 float3314 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6637 float3315 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6638 float3316 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6639 float3317 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7593   word=15   wl=25 address=019f
m6640 LDBL[15] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6641 LDBL[31] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6642 float3318 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6643 float3319 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6644 LDBL[79] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6645 float3320 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6646 float3321 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6647 LDBL[127] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6648 LDBL[143] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6649 float3322 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6650 LDBL[175] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6651 float3323 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6652 LDBL[207] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6653 LDBL[223] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6654 LDBL[239] LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6655 float3324 LDWL[25] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9822   word=0   wl=26 address=01a0
m6656 float3325 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6657 LDBL[16] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6658 float3326 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6659 float3327 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6660 float3328 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6661 LDBL[80] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6662 float3329 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6663 float3330 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6664 float3331 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6665 float3332 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6666 float3333 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6667 LDBL[176] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6668 LDBL[192] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6669 float3334 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6670 float3335 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6671 LDBL[240] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5ef1   word=1   wl=26 address=01a1
m6672 LDBL[1] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6673 float3336 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6674 float3337 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6675 float3338 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6676 LDBL[65] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6677 LDBL[81] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6678 LDBL[97] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6679 LDBL[113] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6680 float3339 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6681 LDBL[145] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6682 LDBL[161] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6683 LDBL[177] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6684 LDBL[193] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6685 float3340 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6686 LDBL[225] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6687 float3341 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=88eb   word=2   wl=26 address=01a2
m6688 LDBL[2] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6689 LDBL[18] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6690 float3342 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6691 LDBL[50] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6692 float3343 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6693 LDBL[82] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6694 LDBL[98] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6695 LDBL[114] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6696 float3344 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6697 float3345 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6698 float3346 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6699 LDBL[178] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6700 float3347 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6701 float3348 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6702 float3349 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6703 LDBL[242] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=bfb8   word=3   wl=26 address=01a3
m6704 float3350 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6705 float3351 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6706 float3352 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6707 LDBL[51] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6708 LDBL[67] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6709 LDBL[83] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6710 float3353 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6711 LDBL[115] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6712 LDBL[131] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6713 LDBL[147] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6714 LDBL[163] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6715 LDBL[179] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6716 LDBL[195] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6717 LDBL[211] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6718 float3354 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6719 LDBL[243] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c2a1   word=4   wl=26 address=01a4
m6720 LDBL[4] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6721 float3355 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6722 float3356 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6723 float3357 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6724 float3358 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6725 LDBL[84] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6726 float3359 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6727 LDBL[116] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6728 float3360 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6729 LDBL[148] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6730 float3361 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6731 float3362 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6732 float3363 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6733 float3364 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6734 LDBL[228] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6735 LDBL[244] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9deb   word=5   wl=26 address=01a5
m6736 LDBL[5] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6737 LDBL[21] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6738 float3365 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6739 LDBL[53] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6740 float3366 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6741 LDBL[85] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6742 LDBL[101] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6743 LDBL[117] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6744 LDBL[133] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6745 float3367 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6746 LDBL[165] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6747 LDBL[181] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6748 LDBL[197] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6749 float3368 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6750 float3369 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6751 LDBL[245] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b9b1   word=6   wl=26 address=01a6
m6752 LDBL[6] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6753 float3370 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6754 float3371 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6755 float3372 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6756 LDBL[70] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6757 LDBL[86] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6758 float3373 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6759 LDBL[118] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6760 LDBL[134] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6761 float3374 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6762 float3375 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6763 LDBL[182] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6764 LDBL[198] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6765 LDBL[214] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6766 float3376 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6767 LDBL[246] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4747   word=7   wl=26 address=01a7
m6768 LDBL[7] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6769 LDBL[23] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6770 LDBL[39] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6771 float3377 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6772 float3378 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6773 float3379 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6774 LDBL[103] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6775 float3380 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6776 LDBL[135] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6777 LDBL[151] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6778 LDBL[167] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6779 float3381 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6780 float3382 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6781 float3383 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6782 LDBL[231] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6783 float3384 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=a4b7   word=8   wl=26 address=01a8
m6784 LDBL[8] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6785 LDBL[24] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6786 LDBL[40] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6787 float3385 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6788 LDBL[72] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6789 LDBL[88] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6790 float3386 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6791 LDBL[120] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6792 float3387 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6793 float3388 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6794 LDBL[168] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6795 float3389 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6796 float3390 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6797 LDBL[216] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6798 float3391 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6799 LDBL[248] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9b39   word=9   wl=26 address=01a9
m6800 LDBL[9] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6801 float3392 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6802 float3393 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6803 LDBL[57] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6804 LDBL[73] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6805 LDBL[89] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6806 float3394 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6807 float3395 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6808 LDBL[137] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6809 LDBL[153] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6810 float3396 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6811 LDBL[185] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6812 LDBL[201] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6813 float3397 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6814 float3398 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6815 LDBL[249] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d6db   word=10   wl=26 address=01aa
m6816 LDBL[10] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6817 LDBL[26] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6818 float3399 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6819 LDBL[58] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6820 LDBL[74] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6821 float3400 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6822 LDBL[106] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6823 LDBL[122] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6824 float3401 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6825 LDBL[154] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6826 LDBL[170] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6827 float3402 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6828 LDBL[202] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6829 float3403 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6830 LDBL[234] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6831 LDBL[250] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fa06   word=11   wl=26 address=01ab
m6832 float3404 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6833 LDBL[27] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6834 LDBL[43] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6835 float3405 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6836 float3406 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6837 float3407 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6838 float3408 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6839 float3409 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6840 float3410 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6841 LDBL[155] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6842 float3411 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6843 LDBL[187] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6844 LDBL[203] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6845 LDBL[219] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6846 LDBL[235] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6847 LDBL[251] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0eb3   word=12   wl=26 address=01ac
m6848 LDBL[12] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6849 LDBL[28] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6850 float3412 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6851 float3413 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6852 LDBL[76] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6853 LDBL[92] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6854 float3414 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6855 LDBL[124] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6856 float3415 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6857 LDBL[156] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6858 LDBL[172] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6859 LDBL[188] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6860 float3416 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6861 float3417 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6862 float3418 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6863 float3419 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=68a9   word=13   wl=26 address=01ad
m6864 LDBL[13] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6865 float3420 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6866 float3421 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6867 LDBL[61] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6868 float3422 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6869 LDBL[93] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6870 float3423 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6871 LDBL[125] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6872 float3424 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6873 float3425 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6874 float3426 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6875 LDBL[189] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6876 float3427 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6877 LDBL[221] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6878 LDBL[237] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6879 float3428 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=479a   word=14   wl=26 address=01ae
m6880 float3429 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6881 LDBL[30] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6882 float3430 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6883 LDBL[62] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6884 LDBL[78] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6885 float3431 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6886 float3432 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6887 LDBL[126] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6888 LDBL[142] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6889 LDBL[158] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6890 LDBL[174] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6891 float3433 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6892 float3434 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6893 float3435 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6894 LDBL[238] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6895 float3436 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=5214   word=15   wl=26 address=01af
m6896 float3437 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6897 float3438 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6898 LDBL[47] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6899 float3439 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6900 LDBL[79] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6901 float3440 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6902 float3441 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6903 float3442 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6904 float3443 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6905 LDBL[159] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6906 float3444 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6907 float3445 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6908 LDBL[207] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6909 float3446 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6910 LDBL[239] LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6911 float3447 LDWL[26] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4668   word=0   wl=27 address=01b0
m6912 float3448 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6913 float3449 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6914 float3450 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6915 LDBL[48] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6916 float3451 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6917 LDBL[80] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6918 LDBL[96] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6919 float3452 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6920 float3453 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6921 LDBL[144] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6922 LDBL[160] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6923 float3454 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6924 float3455 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6925 float3456 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6926 LDBL[224] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6927 float3457 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4af8   word=1   wl=27 address=01b1
m6928 float3458 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6929 float3459 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6930 float3460 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6931 LDBL[49] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6932 LDBL[65] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6933 LDBL[81] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6934 LDBL[97] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6935 LDBL[113] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6936 float3461 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6937 LDBL[145] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6938 float3462 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6939 LDBL[177] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6940 float3463 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6941 float3464 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6942 LDBL[225] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6943 float3465 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8f6a   word=2   wl=27 address=01b2
m6944 float3466 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6945 LDBL[18] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6946 float3467 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6947 LDBL[50] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6948 float3468 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6949 LDBL[82] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6950 LDBL[98] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6951 float3469 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6952 LDBL[130] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6953 LDBL[146] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6954 LDBL[162] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6955 LDBL[178] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6956 float3470 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6957 float3471 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6958 float3472 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6959 LDBL[242] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6414   word=3   wl=27 address=01b3
m6960 float3473 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6961 float3474 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6962 LDBL[35] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6963 float3475 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6964 LDBL[67] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6965 float3476 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6966 float3477 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6967 float3478 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6968 float3479 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6969 float3480 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6970 LDBL[163] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6971 float3481 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6972 float3482 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6973 LDBL[211] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6974 LDBL[227] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6975 float3483 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6c0c   word=4   wl=27 address=01b4
m6976 float3484 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6977 float3485 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6978 LDBL[36] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6979 LDBL[52] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6980 float3486 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6981 float3487 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6982 float3488 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6983 float3489 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6984 float3490 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6985 float3491 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6986 LDBL[164] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6987 LDBL[180] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6988 float3492 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6989 LDBL[212] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6990 LDBL[228] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6991 float3493 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6836   word=5   wl=27 address=01b5
m6992 float3494 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6993 LDBL[21] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6994 LDBL[37] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6995 float3495 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6996 LDBL[69] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6997 LDBL[85] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6998 float3496 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m6999 float3497 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7000 float3498 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7001 float3499 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7002 float3500 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7003 LDBL[181] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7004 float3501 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7005 LDBL[213] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7006 LDBL[229] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7007 float3502 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=dec2   word=6   wl=27 address=01b6
m7008 float3503 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7009 LDBL[22] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7010 float3504 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7011 float3505 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7012 float3506 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7013 float3507 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7014 LDBL[102] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7015 LDBL[118] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7016 float3508 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7017 LDBL[150] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7018 LDBL[166] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7019 LDBL[182] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7020 LDBL[198] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7021 float3509 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7022 LDBL[230] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7023 LDBL[246] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b8e5   word=7   wl=27 address=01b7
m7024 LDBL[7] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7025 float3510 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7026 LDBL[39] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7027 float3511 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7028 float3512 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7029 LDBL[87] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7030 LDBL[103] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7031 LDBL[119] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7032 float3513 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7033 float3514 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7034 float3515 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7035 LDBL[183] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7036 LDBL[199] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7037 LDBL[215] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7038 float3516 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7039 LDBL[247] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8be6   word=8   wl=27 address=01b8
m7040 float3517 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7041 LDBL[24] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7042 LDBL[40] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7043 float3518 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7044 float3519 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7045 LDBL[88] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7046 LDBL[104] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7047 LDBL[120] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7048 LDBL[136] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7049 LDBL[152] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7050 float3520 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7051 LDBL[184] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7052 float3521 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7053 float3522 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7054 float3523 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7055 LDBL[248] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d423   word=9   wl=27 address=01b9
m7056 LDBL[9] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7057 LDBL[25] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7058 float3524 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7059 float3525 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7060 float3526 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7061 LDBL[89] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7062 float3527 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7063 float3528 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7064 float3529 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7065 float3530 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7066 LDBL[169] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7067 float3531 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7068 LDBL[201] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7069 float3532 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7070 LDBL[233] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7071 LDBL[249] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e607   word=10   wl=27 address=01ba
m7072 LDBL[10] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7073 LDBL[26] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7074 LDBL[42] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7075 float3533 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7076 float3534 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7077 float3535 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7078 float3536 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7079 float3537 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7080 float3538 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7081 LDBL[154] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7082 LDBL[170] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7083 float3539 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7084 float3540 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7085 LDBL[218] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7086 LDBL[234] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7087 LDBL[250] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e879   word=11   wl=27 address=01bb
m7088 LDBL[11] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7089 float3541 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7090 float3542 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7091 LDBL[59] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7092 LDBL[75] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7093 LDBL[91] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7094 LDBL[107] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7095 float3543 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7096 float3544 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7097 float3545 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7098 float3546 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7099 LDBL[187] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7100 float3547 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7101 LDBL[219] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7102 LDBL[235] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7103 LDBL[251] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9f88   word=12   wl=27 address=01bc
m7104 float3548 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7105 float3549 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7106 float3550 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7107 LDBL[60] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7108 float3551 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7109 float3552 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7110 float3553 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7111 LDBL[124] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7112 LDBL[140] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7113 LDBL[156] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7114 LDBL[172] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7115 LDBL[188] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7116 LDBL[204] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7117 float3554 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7118 float3555 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7119 LDBL[252] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d70d   word=13   wl=27 address=01bd
m7120 LDBL[13] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7121 float3556 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7122 LDBL[45] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7123 LDBL[61] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7124 float3557 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7125 float3558 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7126 float3559 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7127 float3560 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7128 LDBL[141] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7129 LDBL[157] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7130 LDBL[173] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7131 float3561 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7132 LDBL[205] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7133 float3562 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7134 LDBL[237] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7135 LDBL[253] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3201   word=14   wl=27 address=01be
m7136 LDBL[14] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7137 float3563 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7138 float3564 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7139 float3565 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7140 float3566 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7141 float3567 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7142 float3568 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7143 float3569 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7144 float3570 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7145 LDBL[158] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7146 float3571 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7147 float3572 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7148 LDBL[206] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7149 LDBL[222] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7150 float3573 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7151 float3574 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=cde9   word=15   wl=27 address=01bf
m7152 LDBL[15] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7153 float3575 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7154 float3576 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7155 LDBL[63] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7156 float3577 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7157 LDBL[95] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7158 LDBL[111] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7159 LDBL[127] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7160 LDBL[143] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7161 float3578 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7162 LDBL[175] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7163 LDBL[191] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7164 float3579 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7165 float3580 LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7166 LDBL[239] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7167 LDBL[255] LDWL[27] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4a42   word=0   wl=28 address=01c0
m7168 float3581 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7169 LDBL[16] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7170 float3582 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7171 float3583 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7172 float3584 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7173 float3585 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7174 LDBL[96] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7175 float3586 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7176 float3587 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7177 LDBL[144] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7178 float3588 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7179 LDBL[176] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7180 float3589 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7181 float3590 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7182 LDBL[224] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7183 float3591 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7841   word=1   wl=28 address=01c1
m7184 LDBL[1] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7185 float3592 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7186 float3593 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7187 float3594 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7188 float3595 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7189 float3596 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7190 LDBL[97] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7191 float3597 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7192 float3598 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7193 float3599 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7194 float3600 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7195 LDBL[177] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7196 LDBL[193] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7197 LDBL[209] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7198 LDBL[225] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7199 float3601 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=cc75   word=2   wl=28 address=01c2
m7200 LDBL[2] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7201 float3602 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7202 LDBL[34] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7203 float3603 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7204 LDBL[66] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7205 LDBL[82] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7206 LDBL[98] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7207 float3604 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7208 float3605 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7209 float3606 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7210 LDBL[162] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7211 LDBL[178] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7212 float3607 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7213 float3608 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7214 LDBL[226] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7215 LDBL[242] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=eec8   word=3   wl=28 address=01c3
m7216 float3609 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7217 float3610 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7218 float3611 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7219 LDBL[51] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7220 float3612 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7221 float3613 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7222 LDBL[99] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7223 LDBL[115] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7224 float3614 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7225 LDBL[147] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7226 LDBL[163] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7227 LDBL[179] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7228 float3615 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7229 LDBL[211] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7230 LDBL[227] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7231 LDBL[243] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2549   word=4   wl=28 address=01c4
m7232 LDBL[4] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7233 float3616 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7234 float3617 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7235 LDBL[52] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7236 float3618 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7237 float3619 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7238 LDBL[100] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7239 float3620 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7240 LDBL[132] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7241 float3621 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7242 LDBL[164] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7243 float3622 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7244 float3623 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7245 LDBL[212] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7246 float3624 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7247 float3625 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ac04   word=5   wl=28 address=01c5
m7248 float3626 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7249 float3627 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7250 LDBL[37] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7251 float3628 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7252 float3629 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7253 float3630 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7254 float3631 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7255 float3632 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7256 float3633 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7257 float3634 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7258 LDBL[165] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7259 LDBL[181] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7260 float3635 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7261 LDBL[213] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7262 float3636 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7263 LDBL[245] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=685b   word=6   wl=28 address=01c6
m7264 LDBL[6] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7265 LDBL[22] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7266 float3637 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7267 LDBL[54] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7268 LDBL[70] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7269 float3638 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7270 LDBL[102] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7271 float3639 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7272 float3640 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7273 float3641 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7274 float3642 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7275 LDBL[182] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7276 float3643 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7277 LDBL[214] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7278 LDBL[230] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7279 float3644 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f17f   word=7   wl=28 address=01c7
m7280 LDBL[7] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7281 LDBL[23] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7282 LDBL[39] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7283 LDBL[55] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7284 LDBL[71] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7285 LDBL[87] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7286 LDBL[103] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7287 float3645 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7288 LDBL[135] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7289 float3646 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7290 float3647 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7291 float3648 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7292 LDBL[199] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7293 LDBL[215] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7294 LDBL[231] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7295 LDBL[247] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=95ad   word=8   wl=28 address=01c8
m7296 LDBL[8] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7297 float3649 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7298 LDBL[40] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7299 LDBL[56] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7300 float3650 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7301 LDBL[88] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7302 float3651 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7303 LDBL[120] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7304 LDBL[136] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7305 float3652 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7306 LDBL[168] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7307 float3653 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7308 LDBL[200] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7309 float3654 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7310 float3655 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7311 LDBL[248] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c1dd   word=9   wl=28 address=01c9
m7312 LDBL[9] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7313 float3656 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7314 LDBL[41] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7315 LDBL[57] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7316 LDBL[73] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7317 float3657 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7318 LDBL[105] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7319 LDBL[121] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7320 LDBL[137] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7321 float3658 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7322 float3659 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7323 float3660 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7324 float3661 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7325 float3662 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7326 LDBL[233] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7327 LDBL[249] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=89be   word=10   wl=28 address=01ca
m7328 float3663 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7329 LDBL[26] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7330 LDBL[42] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7331 LDBL[58] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7332 LDBL[74] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7333 LDBL[90] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7334 float3664 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7335 LDBL[122] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7336 LDBL[138] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7337 float3665 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7338 float3666 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7339 LDBL[186] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7340 float3667 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7341 float3668 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7342 float3669 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7343 LDBL[250] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4084   word=11   wl=28 address=01cb
m7344 float3670 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7345 float3671 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7346 LDBL[43] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7347 float3672 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7348 float3673 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7349 float3674 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7350 float3675 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7351 LDBL[123] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7352 float3676 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7353 float3677 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7354 float3678 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7355 float3679 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7356 float3680 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7357 float3681 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7358 LDBL[235] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7359 float3682 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b57d   word=12   wl=28 address=01cc
m7360 LDBL[12] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7361 float3683 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7362 LDBL[44] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7363 LDBL[60] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7364 LDBL[76] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7365 LDBL[92] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7366 LDBL[108] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7367 float3684 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7368 LDBL[140] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7369 float3685 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7370 LDBL[172] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7371 float3686 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7372 LDBL[204] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7373 LDBL[220] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7374 float3687 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7375 LDBL[252] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9718   word=13   wl=28 address=01cd
m7376 float3688 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7377 float3689 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7378 float3690 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7379 LDBL[61] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7380 LDBL[77] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7381 float3691 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7382 float3692 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7383 float3693 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7384 LDBL[141] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7385 LDBL[157] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7386 LDBL[173] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7387 float3694 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7388 LDBL[205] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7389 float3695 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7390 float3696 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7391 LDBL[253] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=16cb   word=14   wl=28 address=01ce
m7392 LDBL[14] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7393 LDBL[30] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7394 float3697 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7395 LDBL[62] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7396 float3698 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7397 float3699 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7398 LDBL[110] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7399 LDBL[126] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7400 float3700 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7401 LDBL[158] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7402 LDBL[174] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7403 float3701 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7404 LDBL[206] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7405 float3702 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7406 float3703 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7407 float3704 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=cafd   word=15   wl=28 address=01cf
m7408 LDBL[15] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7409 float3705 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7410 LDBL[47] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7411 LDBL[63] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7412 LDBL[79] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7413 LDBL[95] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7414 LDBL[111] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7415 LDBL[127] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7416 float3706 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7417 LDBL[159] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7418 float3707 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7419 LDBL[191] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7420 float3708 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7421 float3709 LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7422 LDBL[239] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7423 LDBL[255] LDWL[28] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b86a   word=0   wl=29 address=01d0
m7424 float3710 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7425 LDBL[16] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7426 float3711 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7427 LDBL[48] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7428 float3712 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7429 LDBL[80] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7430 LDBL[96] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7431 float3713 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7432 float3714 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7433 float3715 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7434 float3716 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7435 LDBL[176] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7436 LDBL[192] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7437 LDBL[208] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7438 float3717 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7439 LDBL[240] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=34e6   word=1   wl=29 address=01d1
m7440 float3718 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7441 LDBL[17] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7442 LDBL[33] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7443 float3719 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7444 float3720 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7445 LDBL[81] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7446 LDBL[97] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7447 LDBL[113] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7448 float3721 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7449 float3722 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7450 LDBL[161] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7451 float3723 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7452 LDBL[193] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7453 LDBL[209] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7454 float3724 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7455 float3725 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ff84   word=2   wl=29 address=01d2
m7456 float3726 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7457 float3727 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7458 LDBL[34] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7459 float3728 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7460 float3729 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7461 float3730 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7462 float3731 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7463 LDBL[114] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7464 LDBL[130] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7465 LDBL[146] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7466 LDBL[162] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7467 LDBL[178] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7468 LDBL[194] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7469 LDBL[210] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7470 LDBL[226] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7471 LDBL[242] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6f7f   word=3   wl=29 address=01d3
m7472 LDBL[3] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7473 LDBL[19] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7474 LDBL[35] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7475 LDBL[51] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7476 LDBL[67] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7477 LDBL[83] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7478 LDBL[99] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7479 float3732 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7480 LDBL[131] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7481 LDBL[147] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7482 LDBL[163] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7483 LDBL[179] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7484 float3733 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7485 LDBL[211] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7486 LDBL[227] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7487 float3734 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=64ad   word=4   wl=29 address=01d4
m7488 LDBL[4] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7489 float3735 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7490 LDBL[36] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7491 LDBL[52] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7492 float3736 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7493 LDBL[84] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7494 float3737 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7495 LDBL[116] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7496 float3738 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7497 float3739 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7498 LDBL[164] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7499 float3740 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7500 float3741 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7501 LDBL[212] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7502 LDBL[228] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7503 float3742 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=af4b   word=5   wl=29 address=01d5
m7504 LDBL[5] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7505 LDBL[21] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7506 float3743 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7507 LDBL[53] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7508 float3744 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7509 float3745 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7510 LDBL[101] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7511 float3746 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7512 LDBL[133] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7513 LDBL[149] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7514 LDBL[165] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7515 LDBL[181] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7516 float3747 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7517 LDBL[213] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7518 float3748 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7519 LDBL[245] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=27c2   word=6   wl=29 address=01d6
m7520 float3749 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7521 LDBL[22] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7522 float3750 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7523 float3751 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7524 float3752 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7525 float3753 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7526 LDBL[102] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7527 LDBL[118] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7528 LDBL[134] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7529 LDBL[150] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7530 LDBL[166] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7531 float3754 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7532 float3755 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7533 LDBL[214] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7534 float3756 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7535 float3757 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=644e   word=7   wl=29 address=01d7
m7536 float3758 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7537 LDBL[23] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7538 LDBL[39] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7539 LDBL[55] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7540 float3759 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7541 float3760 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7542 LDBL[103] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7543 float3761 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7544 float3762 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7545 float3763 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7546 LDBL[167] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7547 float3764 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7548 float3765 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7549 LDBL[215] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7550 LDBL[231] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7551 float3766 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9872   word=8   wl=29 address=01d8
m7552 float3767 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7553 LDBL[24] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7554 float3768 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7555 float3769 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7556 LDBL[72] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7557 LDBL[88] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7558 LDBL[104] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7559 float3770 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7560 float3771 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7561 float3772 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7562 float3773 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7563 LDBL[184] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7564 LDBL[200] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7565 float3774 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7566 float3775 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7567 LDBL[248] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=107c   word=9   wl=29 address=01d9
m7568 float3776 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7569 float3777 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7570 LDBL[41] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7571 LDBL[57] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7572 LDBL[73] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7573 LDBL[89] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7574 LDBL[105] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7575 float3778 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7576 float3779 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7577 float3780 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7578 float3781 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7579 float3782 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7580 LDBL[201] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7581 float3783 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7582 float3784 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7583 float3785 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c2bc   word=10   wl=29 address=01da
m7584 float3786 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7585 float3787 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7586 LDBL[42] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7587 LDBL[58] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7588 LDBL[74] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7589 LDBL[90] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7590 float3788 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7591 LDBL[122] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7592 float3789 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7593 LDBL[154] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7594 float3790 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7595 float3791 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7596 float3792 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7597 float3793 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7598 LDBL[234] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7599 LDBL[250] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=0cff   word=11   wl=29 address=01db
m7600 LDBL[11] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7601 LDBL[27] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7602 LDBL[43] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7603 LDBL[59] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7604 LDBL[75] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7605 LDBL[91] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7606 LDBL[107] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7607 LDBL[123] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7608 float3794 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7609 float3795 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7610 LDBL[171] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7611 LDBL[187] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7612 float3796 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7613 float3797 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7614 float3798 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7615 float3799 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=78b5   word=12   wl=29 address=01dc
m7616 LDBL[12] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7617 float3800 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7618 LDBL[44] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7619 float3801 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7620 LDBL[76] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7621 LDBL[92] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7622 float3802 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7623 LDBL[124] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7624 float3803 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7625 float3804 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7626 float3805 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7627 LDBL[188] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7628 LDBL[204] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7629 LDBL[220] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7630 LDBL[236] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7631 float3806 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9a81   word=13   wl=29 address=01dd
m7632 LDBL[13] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7633 float3807 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7634 float3808 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7635 float3809 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7636 float3810 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7637 float3811 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7638 float3812 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7639 LDBL[125] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7640 float3813 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7641 LDBL[157] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7642 float3814 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7643 LDBL[189] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7644 LDBL[205] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7645 float3815 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7646 float3816 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7647 LDBL[253] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=8ec5   word=14   wl=29 address=01de
m7648 LDBL[14] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7649 float3817 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7650 LDBL[46] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7651 float3818 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7652 float3819 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7653 float3820 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7654 LDBL[110] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7655 LDBL[126] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7656 float3821 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7657 LDBL[158] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7658 LDBL[174] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7659 LDBL[190] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7660 float3822 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7661 float3823 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7662 float3824 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7663 LDBL[254] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=b3b1   word=15   wl=29 address=01df
m7664 LDBL[15] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7665 float3825 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7666 float3826 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7667 float3827 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7668 LDBL[79] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7669 LDBL[95] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7670 float3828 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7671 LDBL[127] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7672 LDBL[143] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7673 LDBL[159] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7674 float3829 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7675 float3830 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7676 LDBL[207] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7677 LDBL[223] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7678 float3831 LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7679 LDBL[255] LDWL[29] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e0fc   word=0   wl=30 address=01e0
m7680 float3832 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7681 float3833 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7682 LDBL[32] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7683 LDBL[48] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7684 LDBL[64] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7685 LDBL[80] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7686 LDBL[96] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7687 LDBL[112] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7688 float3834 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7689 float3835 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7690 float3836 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7691 float3837 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7692 float3838 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7693 LDBL[208] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7694 LDBL[224] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7695 LDBL[240] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=63fa   word=1   wl=30 address=01e1
m7696 float3839 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7697 LDBL[17] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7698 float3840 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7699 LDBL[49] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7700 LDBL[65] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7701 LDBL[81] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7702 LDBL[97] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7703 LDBL[113] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7704 LDBL[129] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7705 LDBL[145] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7706 float3841 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7707 float3842 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7708 float3843 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7709 LDBL[209] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7710 LDBL[225] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7711 float3844 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=dc92   word=2   wl=30 address=01e2
m7712 float3845 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7713 LDBL[18] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7714 float3846 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7715 float3847 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7716 LDBL[66] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7717 float3848 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7718 float3849 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7719 LDBL[114] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7720 float3850 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7721 float3851 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7722 LDBL[162] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7723 LDBL[178] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7724 LDBL[194] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7725 float3852 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7726 LDBL[226] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7727 LDBL[242] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=3790   word=3   wl=30 address=01e3
m7728 float3853 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7729 float3854 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7730 float3855 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7731 float3856 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7732 LDBL[67] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7733 float3857 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7734 float3858 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7735 LDBL[115] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7736 LDBL[131] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7737 LDBL[147] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7738 LDBL[163] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7739 float3859 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7740 LDBL[195] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7741 LDBL[211] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7742 float3860 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7743 float3861 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=1e30   word=4   wl=30 address=01e4
m7744 float3862 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7745 float3863 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7746 float3864 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7747 float3865 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7748 LDBL[68] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7749 LDBL[84] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7750 float3866 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7751 float3867 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7752 float3868 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7753 LDBL[148] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7754 LDBL[164] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7755 LDBL[180] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7756 LDBL[196] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7757 float3869 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7758 float3870 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7759 float3871 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e0f1   word=5   wl=30 address=01e5
m7760 LDBL[5] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7761 float3872 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7762 float3873 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7763 float3874 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7764 LDBL[69] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7765 LDBL[85] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7766 LDBL[101] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7767 LDBL[117] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7768 float3875 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7769 float3876 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7770 float3877 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7771 float3878 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7772 float3879 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7773 LDBL[213] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7774 LDBL[229] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7775 LDBL[245] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=43cf   word=6   wl=30 address=01e6
m7776 LDBL[6] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7777 LDBL[22] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7778 LDBL[38] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7779 LDBL[54] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7780 float3880 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7781 float3881 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7782 LDBL[102] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7783 LDBL[118] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7784 LDBL[134] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7785 LDBL[150] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7786 float3882 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7787 float3883 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7788 float3884 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7789 float3885 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7790 LDBL[230] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7791 float3886 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=84b8   word=7   wl=30 address=01e7
m7792 float3887 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7793 float3888 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7794 float3889 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7795 LDBL[55] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7796 LDBL[71] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7797 LDBL[87] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7798 float3890 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7799 LDBL[119] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7800 float3891 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7801 float3892 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7802 LDBL[167] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7803 float3893 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7804 float3894 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7805 float3895 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7806 float3896 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7807 LDBL[247] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2fcc   word=8   wl=30 address=01e8
m7808 float3897 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7809 float3898 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7810 LDBL[40] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7811 LDBL[56] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7812 float3899 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7813 float3900 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7814 LDBL[104] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7815 LDBL[120] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7816 LDBL[136] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7817 LDBL[152] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7818 LDBL[168] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7819 LDBL[184] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7820 float3901 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7821 LDBL[216] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7822 float3902 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7823 float3903 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=f676   word=9   wl=30 address=01e9
m7824 float3904 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7825 LDBL[25] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7826 LDBL[41] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7827 float3905 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7828 LDBL[73] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7829 LDBL[89] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7830 LDBL[105] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7831 float3906 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7832 float3907 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7833 LDBL[153] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7834 LDBL[169] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7835 float3908 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7836 LDBL[201] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7837 LDBL[217] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7838 LDBL[233] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7839 LDBL[249] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6eb0   word=10   wl=30 address=01ea
m7840 float3909 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7841 float3910 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7842 float3911 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7843 float3912 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7844 LDBL[74] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7845 LDBL[90] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7846 float3913 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7847 LDBL[122] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7848 float3914 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7849 LDBL[154] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7850 LDBL[170] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7851 LDBL[186] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7852 float3915 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7853 LDBL[218] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7854 LDBL[234] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7855 float3916 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c3c9   word=11   wl=30 address=01eb
m7856 LDBL[11] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7857 float3917 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7858 float3918 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7859 LDBL[59] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7860 float3919 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7861 float3920 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7862 LDBL[107] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7863 LDBL[123] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7864 LDBL[139] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7865 LDBL[155] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7866 float3921 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7867 float3922 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7868 float3923 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7869 float3924 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7870 LDBL[235] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7871 LDBL[251] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4b0e   word=12   wl=30 address=01ec
m7872 float3925 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7873 LDBL[28] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7874 LDBL[44] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7875 LDBL[60] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7876 float3926 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7877 float3927 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7878 float3928 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7879 float3929 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7880 LDBL[140] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7881 LDBL[156] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7882 float3930 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7883 LDBL[188] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7884 float3931 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7885 float3932 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7886 LDBL[236] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7887 float3933 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7709   word=13   wl=30 address=01ed
m7888 LDBL[13] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7889 float3934 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7890 float3935 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7891 LDBL[61] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7892 float3936 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7893 float3937 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7894 float3938 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7895 float3939 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7896 LDBL[141] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7897 LDBL[157] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7898 LDBL[173] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7899 float3940 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7900 LDBL[205] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7901 LDBL[221] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7902 LDBL[237] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7903 float3941 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=bd22   word=14   wl=30 address=01ee
m7904 float3942 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7905 LDBL[30] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7906 float3943 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7907 float3944 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7908 float3945 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7909 LDBL[94] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7910 float3946 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7911 float3947 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7912 LDBL[142] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7913 float3948 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7914 LDBL[174] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7915 LDBL[190] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7916 LDBL[206] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7917 LDBL[222] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7918 float3949 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7919 LDBL[254] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=7109   word=15   wl=30 address=01ef
m7920 LDBL[15] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7921 float3950 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7922 float3951 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7923 LDBL[63] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7924 float3952 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7925 float3953 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7926 float3954 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7927 float3955 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7928 LDBL[143] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7929 float3956 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7930 float3957 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7931 float3958 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7932 LDBL[207] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7933 LDBL[223] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7934 LDBL[239] LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7935 float3959 LDWL[30] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=d6d3   word=0   wl=31 address=01f0
m7936 LDBL[0] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7937 LDBL[16] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7938 float3960 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7939 float3961 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7940 LDBL[64] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7941 float3962 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7942 LDBL[96] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7943 LDBL[112] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7944 float3963 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7945 LDBL[144] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7946 LDBL[160] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7947 float3964 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7948 LDBL[192] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7949 float3965 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7950 LDBL[224] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7951 LDBL[240] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=830a   word=1   wl=31 address=01f1
m7952 float3966 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7953 LDBL[17] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7954 float3967 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7955 LDBL[49] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7956 float3968 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7957 float3969 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7958 float3970 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7959 float3971 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7960 LDBL[129] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7961 LDBL[145] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7962 float3972 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7963 float3973 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7964 float3974 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7965 float3975 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7966 float3976 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7967 LDBL[241] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=82ce   word=2   wl=31 address=01f2
m7968 float3977 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7969 LDBL[18] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7970 LDBL[34] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7971 LDBL[50] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7972 float3978 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7973 float3979 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7974 LDBL[98] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7975 LDBL[114] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7976 float3980 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7977 LDBL[146] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7978 float3981 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7979 float3982 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7980 float3983 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7981 float3984 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7982 float3985 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7983 LDBL[242] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=4e50   word=3   wl=31 address=01f3
m7984 float3986 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7985 float3987 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7986 float3988 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7987 float3989 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7988 LDBL[67] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7989 float3990 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7990 LDBL[99] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7991 float3991 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7992 float3992 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7993 LDBL[147] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7994 LDBL[163] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7995 LDBL[179] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7996 float3993 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7997 float3994 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7998 LDBL[227] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m7999 float3995 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=9dd0   word=4   wl=31 address=01f4
m8000 float3996 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8001 float3997 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8002 float3998 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8003 float3999 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8004 LDBL[68] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8005 float4000 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8006 LDBL[100] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8007 LDBL[116] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8008 LDBL[132] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8009 float4001 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8010 LDBL[164] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8011 LDBL[180] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8012 LDBL[196] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8013 float4002 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8014 float4003 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8015 LDBL[244] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=fa34   word=5   wl=31 address=01f5
m8016 float4004 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8017 float4005 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8018 LDBL[37] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8019 float4006 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8020 LDBL[69] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8021 LDBL[85] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8022 float4007 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8023 float4008 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8024 float4009 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8025 LDBL[149] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8026 float4010 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8027 LDBL[181] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8028 LDBL[197] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8029 LDBL[213] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8030 LDBL[229] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8031 LDBL[245] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=40c8   word=6   wl=31 address=01f6
m8032 float4011 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8033 float4012 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8034 float4013 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8035 LDBL[54] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8036 float4014 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8037 float4015 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8038 LDBL[102] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8039 LDBL[118] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8040 float4016 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8041 float4017 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8042 float4018 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8043 float4019 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8044 float4020 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8045 float4021 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8046 LDBL[230] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8047 float4022 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=c260   word=7   wl=31 address=01f7
m8048 float4023 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8049 float4024 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8050 float4025 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8051 float4026 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8052 float4027 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8053 LDBL[87] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8054 LDBL[103] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8055 float4028 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8056 float4029 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8057 LDBL[151] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8058 float4030 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8059 float4031 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8060 float4032 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8061 float4033 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8062 LDBL[231] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8063 LDBL[247] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=ebdf   word=8   wl=31 address=01f8
m8064 LDBL[8] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8065 LDBL[24] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8066 LDBL[40] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8067 LDBL[56] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8068 LDBL[72] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8069 float4034 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8070 LDBL[104] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8071 LDBL[120] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8072 LDBL[136] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8073 LDBL[152] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8074 float4035 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8075 LDBL[184] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8076 float4036 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8077 LDBL[216] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8078 LDBL[232] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8079 LDBL[248] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=2611   word=9   wl=31 address=01f9
m8080 LDBL[9] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8081 float4037 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8082 float4038 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8083 float4039 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8084 LDBL[73] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8085 float4040 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8086 float4041 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8087 float4042 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8088 float4043 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8089 LDBL[153] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8090 LDBL[169] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8091 float4044 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8092 float4045 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8093 LDBL[217] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8094 float4046 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8095 float4047 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=af0e   word=10   wl=31 address=01fa
m8096 float4048 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8097 LDBL[26] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8098 LDBL[42] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8099 LDBL[58] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8100 float4049 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8101 float4050 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8102 float4051 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8103 float4052 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8104 LDBL[138] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8105 LDBL[154] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8106 LDBL[170] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8107 LDBL[186] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8108 float4053 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8109 LDBL[218] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8110 float4054 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8111 LDBL[250] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=e6b1   word=11   wl=31 address=01fb
m8112 LDBL[11] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8113 float4055 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8114 float4056 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8115 float4057 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8116 LDBL[75] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8117 LDBL[91] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8118 float4058 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8119 LDBL[123] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8120 float4059 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8121 LDBL[155] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8122 LDBL[171] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8123 float4060 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8124 float4061 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8125 LDBL[219] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8126 LDBL[235] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8127 LDBL[251] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=6430   word=12   wl=31 address=01fc
m8128 float4062 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8129 float4063 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8130 float4064 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8131 float4065 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8132 LDBL[76] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8133 LDBL[92] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8134 float4066 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8135 float4067 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8136 float4068 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8137 float4069 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8138 LDBL[172] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8139 float4070 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8140 float4071 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8141 LDBL[220] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8142 LDBL[236] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8143 float4072 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=841f   word=13   wl=31 address=01fd
m8144 LDBL[13] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8145 LDBL[29] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8146 LDBL[45] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8147 LDBL[61] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8148 LDBL[77] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8149 float4073 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8150 float4074 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8151 float4075 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8152 float4076 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8153 float4077 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8154 LDBL[173] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8155 float4078 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8156 float4079 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8157 float4080 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8158 float4081 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8159 LDBL[253] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=388c   word=14   wl=31 address=01fe
m8160 float4082 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8161 float4083 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8162 LDBL[46] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8163 LDBL[62] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8164 float4084 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8165 float4085 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8166 float4086 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8167 LDBL[126] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8168 float4087 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8169 float4088 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8170 float4089 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8171 LDBL[190] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8172 LDBL[206] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8173 LDBL[222] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8174 float4090 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8175 float4091 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
*   pattern=47e6   word=15   wl=31 address=01ff
m8176 float4092 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8177 LDBL[31] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8178 LDBL[47] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8179 float4093 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8180 float4094 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8181 LDBL[95] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8182 LDBL[111] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8183 LDBL[127] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8184 LDBL[143] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8185 LDBL[159] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8186 LDBL[175] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8187 float4095 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8188 float4096 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8189 float4097 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8190 LDBL[239] LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
m8191 float4098 LDWL[31] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=1
Vkeep1 LDWL[32] 0 0
*   pattern=5c81   word=0   wl=32 address=0200
m8192 LDBL[0] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8193 LDBL[16] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8194 LDBL[32] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8195 LDBL[48] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8196 LDBL[64] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8197 LDBL[80] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8198 LDBL[96] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8199 LDBL[112] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8200 LDBL[128] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8201 LDBL[144] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8202 LDBL[160] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8203 LDBL[176] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8204 LDBL[192] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8205 LDBL[208] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8206 LDBL[224] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8207 LDBL[240] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=8998   word=1   wl=32 address=0201
m8208 LDBL[1] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8209 LDBL[17] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8210 LDBL[33] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8211 LDBL[49] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8212 LDBL[65] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8213 LDBL[81] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8214 LDBL[97] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8215 LDBL[113] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8216 LDBL[129] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8217 LDBL[145] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8218 LDBL[161] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8219 LDBL[177] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8220 LDBL[193] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8221 LDBL[209] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8222 LDBL[225] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8223 LDBL[241] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=71b0   word=2   wl=32 address=0202
m8224 LDBL[2] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8225 LDBL[18] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8226 LDBL[34] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8227 LDBL[50] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8228 LDBL[66] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8229 LDBL[82] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8230 LDBL[98] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8231 LDBL[114] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8232 LDBL[130] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8233 LDBL[146] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8234 LDBL[162] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8235 LDBL[178] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8236 LDBL[194] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8237 LDBL[210] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8238 LDBL[226] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8239 LDBL[242] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=717e   word=3   wl=32 address=0203
m8240 LDBL[3] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8241 LDBL[19] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8242 LDBL[35] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8243 LDBL[51] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8244 LDBL[67] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8245 LDBL[83] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8246 LDBL[99] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8247 LDBL[115] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8248 LDBL[131] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8249 LDBL[147] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8250 LDBL[163] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8251 LDBL[179] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8252 LDBL[195] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8253 LDBL[211] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8254 LDBL[227] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8255 LDBL[243] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=70ce   word=4   wl=32 address=0204
m8256 LDBL[4] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8257 LDBL[20] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8258 LDBL[36] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8259 LDBL[52] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8260 LDBL[68] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8261 LDBL[84] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8262 LDBL[100] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8263 LDBL[116] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8264 LDBL[132] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8265 LDBL[148] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8266 LDBL[164] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8267 LDBL[180] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8268 LDBL[196] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8269 LDBL[212] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8270 LDBL[228] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8271 LDBL[244] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=b1d5   word=5   wl=32 address=0205
m8272 LDBL[5] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8273 LDBL[21] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8274 LDBL[37] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8275 LDBL[53] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8276 LDBL[69] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8277 LDBL[85] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8278 LDBL[101] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8279 LDBL[117] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8280 LDBL[133] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8281 LDBL[149] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8282 LDBL[165] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8283 LDBL[181] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8284 LDBL[197] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8285 LDBL[213] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8286 LDBL[229] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8287 LDBL[245] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=bfb2   word=6   wl=32 address=0206
m8288 LDBL[6] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8289 LDBL[22] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8290 LDBL[38] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8291 LDBL[54] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8292 LDBL[70] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8293 LDBL[86] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8294 LDBL[102] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8295 LDBL[118] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8296 LDBL[134] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8297 LDBL[150] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8298 LDBL[166] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8299 LDBL[182] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8300 LDBL[198] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8301 LDBL[214] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8302 LDBL[230] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8303 LDBL[246] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=afe4   word=7   wl=32 address=0207
m8304 LDBL[7] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8305 LDBL[23] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8306 LDBL[39] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8307 LDBL[55] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8308 LDBL[71] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8309 LDBL[87] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8310 LDBL[103] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8311 LDBL[119] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8312 LDBL[135] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8313 LDBL[151] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8314 LDBL[167] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8315 LDBL[183] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8316 LDBL[199] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8317 LDBL[215] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8318 LDBL[231] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8319 LDBL[247] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=6f1c   word=8   wl=32 address=0208
m8320 LDBL[8] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8321 LDBL[24] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8322 LDBL[40] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8323 LDBL[56] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8324 LDBL[72] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8325 LDBL[88] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8326 LDBL[104] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8327 LDBL[120] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8328 LDBL[136] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8329 LDBL[152] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8330 LDBL[168] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8331 LDBL[184] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8332 LDBL[200] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8333 LDBL[216] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8334 LDBL[232] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8335 LDBL[248] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=17fc   word=9   wl=32 address=0209
m8336 LDBL[9] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8337 LDBL[25] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8338 LDBL[41] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8339 LDBL[57] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8340 LDBL[73] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8341 LDBL[89] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8342 LDBL[105] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8343 LDBL[121] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8344 LDBL[137] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8345 LDBL[153] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8346 LDBL[169] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8347 LDBL[185] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8348 LDBL[201] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8349 LDBL[217] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8350 LDBL[233] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8351 LDBL[249] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=8ba0   word=10   wl=32 address=020a
m8352 LDBL[10] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8353 LDBL[26] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8354 LDBL[42] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8355 LDBL[58] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8356 LDBL[74] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8357 LDBL[90] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8358 LDBL[106] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8359 LDBL[122] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8360 LDBL[138] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8361 LDBL[154] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8362 LDBL[170] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8363 LDBL[186] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8364 LDBL[202] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8365 LDBL[218] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8366 LDBL[234] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8367 LDBL[250] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=7ad4   word=11   wl=32 address=020b
m8368 LDBL[11] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8369 LDBL[27] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8370 LDBL[43] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8371 LDBL[59] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8372 LDBL[75] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8373 LDBL[91] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8374 LDBL[107] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8375 LDBL[123] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8376 LDBL[139] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8377 LDBL[155] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8378 LDBL[171] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8379 LDBL[187] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8380 LDBL[203] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8381 LDBL[219] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8382 LDBL[235] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8383 LDBL[251] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=add2   word=12   wl=32 address=020c
m8384 LDBL[12] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8385 LDBL[28] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8386 LDBL[44] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8387 LDBL[60] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8388 LDBL[76] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8389 LDBL[92] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8390 LDBL[108] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8391 LDBL[124] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8392 LDBL[140] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8393 LDBL[156] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8394 LDBL[172] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8395 LDBL[188] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8396 LDBL[204] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8397 LDBL[220] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8398 LDBL[236] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8399 LDBL[252] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=7501   word=13   wl=32 address=020d
m8400 LDBL[13] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8401 LDBL[29] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8402 LDBL[45] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8403 LDBL[61] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8404 LDBL[77] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8405 LDBL[93] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8406 LDBL[109] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8407 LDBL[125] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8408 LDBL[141] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8409 LDBL[157] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8410 LDBL[173] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8411 LDBL[189] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8412 LDBL[205] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8413 LDBL[221] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8414 LDBL[237] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8415 LDBL[253] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=bb54   word=14   wl=32 address=020e
m8416 LDBL[14] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8417 LDBL[30] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8418 LDBL[46] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8419 LDBL[62] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8420 LDBL[78] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8421 LDBL[94] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8422 LDBL[110] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8423 LDBL[126] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8424 LDBL[142] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8425 LDBL[158] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8426 LDBL[174] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8427 LDBL[190] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8428 LDBL[206] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8429 LDBL[222] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8430 LDBL[238] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8431 LDBL[254] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
*   pattern=9942   word=15   wl=32 address=020f
m8432 LDBL[15] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8433 LDBL[31] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8434 LDBL[47] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8435 LDBL[63] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8436 LDBL[79] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8437 LDBL[95] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8438 LDBL[111] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8439 LDBL[127] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8440 LDBL[143] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8441 LDBL[159] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8442 LDBL[175] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8443 LDBL[191] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8444 LDBL[207] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8445 LDBL[223] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8446 LDBL[239] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480
m8447 LDBL[255] LDWL[32] 0 0 cmosn AD=17.6e-12 AS=17.6e-12 L=2.4e-06 PD=16.8e-06 PS=16.8e-06 W=4e-06
+ m=480

**** end user architecture code
.ends


* expanding   symbol:  lvnot.sym # of pins=2
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/lvnot.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/lvnot.sch
.subckt lvnot  y a  VCCPIN  VSSPIN      wn=10u lln=1.2u wp=10u lp=1.2u
*.opin y
*.ipin a
m2 y a VCCPIN VCCPIN cmosp w=wp l=lp ad='wp *4.6u' as='wp *4.6u' pd='wp *2+9.2u' ps='wp *2+9.2u' m=1
m1 y a VSSPIN VSSPIN cmosn w=wn l=lln ad='wn *4.3u' as='wn *4.3u' pd='wn *2+8.6u' ps='wn *2+8.6u' m=1
.ends


* expanding   symbol:  bts.sym # of pins=3
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/bts.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/bts.sch
.subckt bts  Z A E  VCCPIN  VSSPIN
*.ipin A
*.ipin E
*.opin Z
m7 NN EN PP VCCPIN cmosp w=56u l=2.4u ad='56u *2.2u' as='56u *2.2u' pd='56u *2+4.4u' ps='56u *2+4.4u'
+ m=1
m8 PP A VCCPIN VCCPIN cmosp w=56u l=2.4u ad='56u *2.2u' as='56u *2.2u' pd='56u *2+4.4u' ps='56u *2+4.4u'
+ m=1
m9 NN A VSSPIN 0 cmosn w=20u l=2.4u ad='20u *4.4u' as='20u *4.4u' pd='20u *2 + 8.8u' ps='20u *2 + 8.8u'
+ m=1
m1 PP E NN 0 cmosn w=24u l=2.4u ad='24u *4.4u' as='24u *4.4u' pd='24u *2 + 8.8u' ps='24u *2 + 8.8u' m=1
m11 Z PP VCCPIN VCCPIN cmosp w=200u l=2.4u ad='200u *2.2u' as='200u *2.2u' pd='200u *2+4.4u' ps='200u *2+4.4u'
+ m=1
m12 Z NN VSSPIN 0 cmosn w=80u l=2.4u ad='80u *4.4u' as='80u *4.4u' pd='80u *2 + 8.8u' ps='80u *2 + 8.8u'
+ m=1
m13 NN EN VSSPIN 0 cmosn w=20u l=2.4u ad='20u *4.4u' as='20u *4.4u' pd='20u *2 + 8.8u' ps='20u *2 + 8.8u'
+ m=1
m14 PP E VCCPIN VCCPIN cmosp w=50u l=2.4u ad='50u *2.2u' as='50u *2.2u' pd='50u *2+4.4u' ps='50u *2+4.4u'
+ m=1
m15 EN E VCCPIN VCCPIN cmosp w=50u l=2.4u ad='50u *2.2u' as='50u *2.2u' pd='50u *2+4.4u' ps='50u *2+4.4u'
+ m=1
m16 EN E VSSPIN 0 cmosn w=20u l=2.4u ad='20u *4.4u' as='20u *4.4u' pd='20u *2 + 8.8u' ps='20u *2 + 8.8u'
+ m=1
c0 E VSSPIN 3f m=1
c4 NN VSSPIN 3f m=1
c5 PP VSSPIN 3f m=1
c6 EN VSSPIN 3f m=1
.ends


* expanding   symbol:  passhs.sym # of pins=4
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/passhs.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/passhs.sch
.subckt passhs  Z A EN E  VCCPIN  VSSPIN   WN=2u LN=1.2u WP=2u LP=1.2u
*.iopin Z
*.iopin A
*.ipin EN
*.ipin E
m60 Z EN A VCCPIN cmosp w=WP l=2.4u ad='WP *4.6u' as='WP *4.6u' pd='WP *2+9.2u' ps='WP *2+9.2u' m=1
m1 A E Z VSSPIN cmosn w=WN l=2.4u ad='WN *4.3u' as='WN *4.3u' pd='WN *2+8.6u' ps='WN *2+8.6u' m=1
.ends


* expanding   symbol:  rom2_sacell.sym # of pins=7
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_sacell.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/rom2_sacell.sch
.subckt rom2_sacell  LDRESET LDPRECH VCC VSS LDQI LDQ_B LDYMS
*.ipin LDRESET
*.ipin LDPRECH
*.ipin VCC
*.ipin VSS
*.opin LDQI
*.opin LDQ_B
*.iopin LDYMS
m3 VCC LDPRECH LDYMS VSS cmosn w=WPRECH l=2u ad='WPRECH *4.3u' as='WPRECH *4.3u' pd='WPRECH *2+8.6u'
+ ps='WPRECH *2+8.6u' m=10
m1 LDQI VCC LDYMS VSS cmosn w=WPRECH l=2u ad='WPRECH *4.3u' as='WPRECH *4.3u' pd='WPRECH *2+8.6u' ps='WPRECH *2+8.6u'
+ m=2
m5 LDQI LDRESET VCC VCC cmosp w=6.6u l=8.8u ad='6.6u *4.4u' as='6.6u *4.4u' pd='6.6u *2 + 8.8u' ps='6.6u *2 + 8.8u'
+ m=1
m11 LDYMS LDRESET VSS 0 cmosn w=16u l=2.4u ad='16u *4.4u' as='16u *4.4u' pd='16u *2 + 8.8u' ps='16u *2 + 8.8u'
+ m=1
c2 LDQI VSS 3f m=1
m2 LDQ_B LDQI VSS 0 cmosn w=8u l=2.4u ad='8u *4.4u' as='8u *4.4u' pd='8u *2 + 8.8u' ps='8u *2 + 8.8u'
+ m=1
m4 LDQ_B LDQI VCC VCC cmosp w=40u l=2.4u ad='40u *4.6u' as='40u *4.6u' pd='40u *2+9.2u' ps='40u *2+9.2u'
+ m=1
.ends


* expanding   symbol:  LD2QHDX4stef.sym # of pins=8
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/LD2QHDX4stef.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/LD2QHDX4stef.sch
.subckt LD2QHDX4stef  D G CD Q vcc vss vccsup vsssup
*.ipin D
*.ipin G
*.ipin CD
*.opin Q
*.iopin vcc
*.iopin vss
*.iopin vccsup
*.iopin vsssup
c2 BN vss 3f m=1
c3 DDN vss 5f m=1
c5 GN vss 5f m=1
c7 FN vss 3f m=1
x8 DDN BN G GN vccsup vsssup passhs WN=12u LN=1.2u WP=12u LP=1.2u
m17 DDN D net2 vsssup cmosn w=8.4u l=2.4u ad='8.4u *2.2u' as='8.4u *2.2u' pd='8.4u *2+4.4u' ps='8.4u *2+4.4u'
+ m=1
m1 DDN D net3 vccsup cmosp w=20u l=2.4u ad='20u *2.2u' as='20u *2.2u' pd='20u *2+4.4u' ps='20u *2+4.4u'
+ m=1
m2 net2 G net1 vsssup cmosn w=8.4u l=2.4u ad='8.4u *2.2u' as='8.4u *2.2u' pd='8.4u *2+4.4u' ps='8.4u *2+4.4u'
+ m=1
m3 net3 GN vcc vccsup cmosp w=20u l=2.4u ad='20u *2.2u' as='20u *2.2u' pd='20u *2+4.4u' ps='20u *2+4.4u'
+ m=1
m4 BN FN net1 vsssup cmosn w=8.4u l=2.4u ad='8.4u *2.2u' as='8.4u *2.2u' pd='8.4u *2+4.4u' ps='8.4u *2+4.4u'
+ m=1
m5 BN FN vcc vccsup cmosp w=8.4u l=2.4u ad='8.4u *2.2u' as='8.4u *2.2u' pd='8.4u *2+4.4u' ps='8.4u *2+4.4u'
+ m=1
m8 net1 CD vss vsssup cmosn w=24u l=2.4u ad='24u *2.2u' as='24u *2.2u' pd='24u *2+4.4u' ps='24u *2+4.4u'
+ m=1
m11 DDN CD vcc vccsup cmosp w=8.4u l=2.4u ad='8.4u *2.2u' as='8.4u *2.2u' pd='8.4u *2+4.4u' ps='8.4u *2+4.4u'
+ m=1
x10 FN DDN vcc vss lvnot wn=8.4u lln=2.4u wp=8.4u lp=2.4u m=1
x1 GN G vcc vss lvnot wn=40u lln=2.4u wp=40u lp=2.4u m=1
x2 Q DDN vcc vss lvnot wn=40u lln=2.4u wp=100u lp=2.4u m=1
.save  v(ddn)
.save  v(fn)
.ends


* expanding   symbol:  lvnand2.sym # of pins=3
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/lvnand2.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/lvnand2.sch
.subckt lvnand2  y a b  VCCPIN  VSSPIN      wna=8u lna=1.2u wpa=10u lpa=1.2u  wnb=8u lnb=1.2u
+ wpb=10u lpb=1.2u
*.opin y
*.ipin a
*.ipin b
m2 y a VCCPIN VCCPIN cmosp w=wpa l=lpa ad='wpa *4.6u' as='wpa *4.6u' pd='wpa *2+9.2u' ps='wpa *2+9.2u'
+ m=1
m1 y b VCCPIN VCCPIN cmosp w=wpb l=lpb ad='wpb *4.6u' as='wpb *4.6u' pd='wpb *2+9.2u' ps='wpb *2+9.2u'
+ m=1
m3 y a net1 VSSPIN cmosn w=wna l=lna ad='wna *4.3u' as='wna *4.3u' pd='wna *2+8.6u' ps='wna *2+8.6u'
+ m=1
m4 net1 b VSSPIN VSSPIN cmosn w=wnb l=lnb ad='wnb *4.3u' as='wnb *4.3u' pd='wnb *2+8.6u' ps='wnb *2+8.6u'
+ m=1
.ends


* expanding   symbol:  lvnor2.sym # of pins=3
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/lvnor2.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/lvnor2.sch
.subckt lvnor2  y a b  VCCPIN  VSSPIN      wna=2u lna=1.2u wpa=6u lpa=1.2u  wnb=2u lnb=1.2u wpb=6u
+ lpb=1.2u
*.opin y
*.ipin a
*.ipin b
m2 net1 a VCCPIN VCCPIN cmosp w=wpa l=lpa ad='wpa *2.2u' as='wpa *2.2u' pd='wpa *2+4.4u' ps='wpa *2+4.4u'
+ m=1
m1 y b net1 VCCPIN cmosp w=wpb l=lpb ad='wpb *2.2u' as='wpb *2.2u' pd='wpb *2+4.4u' ps='wpb *2+4.4u'
+ m=1
m3 y a VSSPIN VSSPIN cmosn w=wna l=lna ad='wna *2.2u' as='wna *2.2u' pd='wna *2+4.4u' ps='wna *2+4.4u'
+ m=1
m4 y b VSSPIN VSSPIN cmosn w=wnb l=lnb ad='wnb *2.2u' as='wnb *2.2u' pd='wnb *2+4.4u' ps='wnb *2+4.4u'
+ m=1
.ends


* expanding   symbol:  lvnand3.sym # of pins=4
** sym_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/lvnand3.sym
** sch_path:
*+ /foss/tools/xschem/1cb9645e9f84d2dfcb3aecc6e0414d4dede32529/share/doc/xschem/rom8k/lvnand3.sch
.subckt lvnand3  y a b c  VCCPIN  VSSPIN      wn=18u lln=1.2u wp=10u lp=1.2u
*.opin y
*.ipin a
*.ipin b
*.ipin c
m1 net2 a VSSPIN VSSPIN cmosn w=wn l=lln ad='wn *2.2u' as='wn *2.2u' pd='wn *2+4.4u' ps='wn *2+4.4u'
+ m=1
m2 y a VCCPIN VCCPIN cmosp w=wp l=lp ad='wp *2.2u' as='wp *2.2u' pd='wp *2+4.4u' ps='wp *2+4.4u' m=1
m3 y b VCCPIN VCCPIN cmosp w=wp l=lp ad='wp *2.2u' as='wp *2.2u' pd='wp *2+4.4u' ps='wp *2+4.4u' m=1
m5 y c net1 VSSPIN cmosn w=wn l=lln ad='wn *2.2u' as='wn *2.2u' pd='wn *2+4.4u' ps='wn *2+4.4u' m=1
m4 y c VCCPIN VCCPIN cmosp w=wp l=lp ad='wp *2.2u' as='wp *2.2u' pd='wp *2+4.4u' ps='wp *2+4.4u' m=1
m6 net1 b net2 VSSPIN cmosn w=wn l=lln ad='wn *2.2u' as='wn *2.2u' pd='wn *2+4.4u' ps='wn *2+4.4u' m=1
.ends

.end
