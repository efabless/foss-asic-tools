magic
tech sky130A
magscale 1 2
timestamp 1620937039
<< error_p >>
rect -29 581 29 587
rect -29 547 -17 581
rect -29 541 29 547
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect -29 -587 29 -581
<< nwell >>
rect -144 -600 144 600
<< pmoshvt >>
rect -50 -500 50 500
<< pdiff >>
rect -108 488 -50 500
rect -108 -488 -96 488
rect -62 -488 -50 488
rect -108 -500 -50 -488
rect 50 488 108 500
rect 50 -488 62 488
rect 96 -488 108 488
rect 50 -500 108 -488
<< pdiffc >>
rect -96 -488 -62 488
rect 62 -488 96 488
<< poly >>
rect -36 581 36 597
rect -36 564 -20 581
rect -50 547 -20 564
rect 20 564 36 581
rect 20 547 50 564
rect -50 500 50 547
rect -50 -547 50 -500
rect -50 -564 -20 -547
rect -36 -581 -20 -564
rect 20 -564 50 -547
rect 20 -581 36 -564
rect -36 -597 36 -581
<< polycont >>
rect -20 547 20 581
rect -20 -581 20 -547
<< locali >>
rect -36 547 -20 581
rect 20 547 36 581
rect -96 488 -62 504
rect -96 -504 -62 -488
rect 62 488 96 504
rect 62 -504 96 -488
rect -36 -581 -20 -547
rect 20 -581 36 -547
<< viali >>
rect -17 547 17 581
rect -96 -488 -62 488
rect 62 -488 96 488
rect -17 -581 17 -547
<< metal1 >>
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect -102 488 -56 500
rect -102 -488 -96 488
rect -62 -488 -56 488
rect -102 -500 -56 -488
rect 56 488 102 500
rect 56 -488 62 488
rect 96 -488 102 488
rect 56 -500 102 -488
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_hvt
string parameters w 5 l 0.5 m 1 nf 1 diffcov 100 polycov 60 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
