magic
tech sky130A
magscale 1 2
timestamp 1621729938
<< mvnmos >>
rect -6923 -700 -6823 700
rect -6765 -700 -6665 700
rect -6607 -700 -6507 700
rect -6449 -700 -6349 700
rect -6291 -700 -6191 700
rect -6133 -700 -6033 700
rect -5975 -700 -5875 700
rect -5817 -700 -5717 700
rect -5659 -700 -5559 700
rect -5501 -700 -5401 700
rect -5343 -700 -5243 700
rect -5185 -700 -5085 700
rect -5027 -700 -4927 700
rect -4869 -700 -4769 700
rect -4711 -700 -4611 700
rect -4553 -700 -4453 700
rect -4395 -700 -4295 700
rect -4237 -700 -4137 700
rect -4079 -700 -3979 700
rect -3921 -700 -3821 700
rect -3763 -700 -3663 700
rect -3605 -700 -3505 700
rect -3447 -700 -3347 700
rect -3289 -700 -3189 700
rect -3131 -700 -3031 700
rect -2973 -700 -2873 700
rect -2815 -700 -2715 700
rect -2657 -700 -2557 700
rect -2499 -700 -2399 700
rect -2341 -700 -2241 700
rect -2183 -700 -2083 700
rect -2025 -700 -1925 700
rect -1867 -700 -1767 700
rect -1709 -700 -1609 700
rect -1551 -700 -1451 700
rect -1393 -700 -1293 700
rect -1235 -700 -1135 700
rect -1077 -700 -977 700
rect -919 -700 -819 700
rect -761 -700 -661 700
rect -603 -700 -503 700
rect -445 -700 -345 700
rect -287 -700 -187 700
rect -129 -700 -29 700
rect 29 -700 129 700
rect 187 -700 287 700
rect 345 -700 445 700
rect 503 -700 603 700
rect 661 -700 761 700
rect 819 -700 919 700
rect 977 -700 1077 700
rect 1135 -700 1235 700
rect 1293 -700 1393 700
rect 1451 -700 1551 700
rect 1609 -700 1709 700
rect 1767 -700 1867 700
rect 1925 -700 2025 700
rect 2083 -700 2183 700
rect 2241 -700 2341 700
rect 2399 -700 2499 700
rect 2557 -700 2657 700
rect 2715 -700 2815 700
rect 2873 -700 2973 700
rect 3031 -700 3131 700
rect 3189 -700 3289 700
rect 3347 -700 3447 700
rect 3505 -700 3605 700
rect 3663 -700 3763 700
rect 3821 -700 3921 700
rect 3979 -700 4079 700
rect 4137 -700 4237 700
rect 4295 -700 4395 700
rect 4453 -700 4553 700
rect 4611 -700 4711 700
rect 4769 -700 4869 700
rect 4927 -700 5027 700
rect 5085 -700 5185 700
rect 5243 -700 5343 700
rect 5401 -700 5501 700
rect 5559 -700 5659 700
rect 5717 -700 5817 700
rect 5875 -700 5975 700
rect 6033 -700 6133 700
rect 6191 -700 6291 700
rect 6349 -700 6449 700
rect 6507 -700 6607 700
rect 6665 -700 6765 700
rect 6823 -700 6923 700
<< mvndiff >>
rect -6981 688 -6923 700
rect -6981 -688 -6969 688
rect -6935 -688 -6923 688
rect -6981 -700 -6923 -688
rect -6823 688 -6765 700
rect -6823 -688 -6811 688
rect -6777 -688 -6765 688
rect -6823 -700 -6765 -688
rect -6665 688 -6607 700
rect -6665 -688 -6653 688
rect -6619 -688 -6607 688
rect -6665 -700 -6607 -688
rect -6507 688 -6449 700
rect -6507 -688 -6495 688
rect -6461 -688 -6449 688
rect -6507 -700 -6449 -688
rect -6349 688 -6291 700
rect -6349 -688 -6337 688
rect -6303 -688 -6291 688
rect -6349 -700 -6291 -688
rect -6191 688 -6133 700
rect -6191 -688 -6179 688
rect -6145 -688 -6133 688
rect -6191 -700 -6133 -688
rect -6033 688 -5975 700
rect -6033 -688 -6021 688
rect -5987 -688 -5975 688
rect -6033 -700 -5975 -688
rect -5875 688 -5817 700
rect -5875 -688 -5863 688
rect -5829 -688 -5817 688
rect -5875 -700 -5817 -688
rect -5717 688 -5659 700
rect -5717 -688 -5705 688
rect -5671 -688 -5659 688
rect -5717 -700 -5659 -688
rect -5559 688 -5501 700
rect -5559 -688 -5547 688
rect -5513 -688 -5501 688
rect -5559 -700 -5501 -688
rect -5401 688 -5343 700
rect -5401 -688 -5389 688
rect -5355 -688 -5343 688
rect -5401 -700 -5343 -688
rect -5243 688 -5185 700
rect -5243 -688 -5231 688
rect -5197 -688 -5185 688
rect -5243 -700 -5185 -688
rect -5085 688 -5027 700
rect -5085 -688 -5073 688
rect -5039 -688 -5027 688
rect -5085 -700 -5027 -688
rect -4927 688 -4869 700
rect -4927 -688 -4915 688
rect -4881 -688 -4869 688
rect -4927 -700 -4869 -688
rect -4769 688 -4711 700
rect -4769 -688 -4757 688
rect -4723 -688 -4711 688
rect -4769 -700 -4711 -688
rect -4611 688 -4553 700
rect -4611 -688 -4599 688
rect -4565 -688 -4553 688
rect -4611 -700 -4553 -688
rect -4453 688 -4395 700
rect -4453 -688 -4441 688
rect -4407 -688 -4395 688
rect -4453 -700 -4395 -688
rect -4295 688 -4237 700
rect -4295 -688 -4283 688
rect -4249 -688 -4237 688
rect -4295 -700 -4237 -688
rect -4137 688 -4079 700
rect -4137 -688 -4125 688
rect -4091 -688 -4079 688
rect -4137 -700 -4079 -688
rect -3979 688 -3921 700
rect -3979 -688 -3967 688
rect -3933 -688 -3921 688
rect -3979 -700 -3921 -688
rect -3821 688 -3763 700
rect -3821 -688 -3809 688
rect -3775 -688 -3763 688
rect -3821 -700 -3763 -688
rect -3663 688 -3605 700
rect -3663 -688 -3651 688
rect -3617 -688 -3605 688
rect -3663 -700 -3605 -688
rect -3505 688 -3447 700
rect -3505 -688 -3493 688
rect -3459 -688 -3447 688
rect -3505 -700 -3447 -688
rect -3347 688 -3289 700
rect -3347 -688 -3335 688
rect -3301 -688 -3289 688
rect -3347 -700 -3289 -688
rect -3189 688 -3131 700
rect -3189 -688 -3177 688
rect -3143 -688 -3131 688
rect -3189 -700 -3131 -688
rect -3031 688 -2973 700
rect -3031 -688 -3019 688
rect -2985 -688 -2973 688
rect -3031 -700 -2973 -688
rect -2873 688 -2815 700
rect -2873 -688 -2861 688
rect -2827 -688 -2815 688
rect -2873 -700 -2815 -688
rect -2715 688 -2657 700
rect -2715 -688 -2703 688
rect -2669 -688 -2657 688
rect -2715 -700 -2657 -688
rect -2557 688 -2499 700
rect -2557 -688 -2545 688
rect -2511 -688 -2499 688
rect -2557 -700 -2499 -688
rect -2399 688 -2341 700
rect -2399 -688 -2387 688
rect -2353 -688 -2341 688
rect -2399 -700 -2341 -688
rect -2241 688 -2183 700
rect -2241 -688 -2229 688
rect -2195 -688 -2183 688
rect -2241 -700 -2183 -688
rect -2083 688 -2025 700
rect -2083 -688 -2071 688
rect -2037 -688 -2025 688
rect -2083 -700 -2025 -688
rect -1925 688 -1867 700
rect -1925 -688 -1913 688
rect -1879 -688 -1867 688
rect -1925 -700 -1867 -688
rect -1767 688 -1709 700
rect -1767 -688 -1755 688
rect -1721 -688 -1709 688
rect -1767 -700 -1709 -688
rect -1609 688 -1551 700
rect -1609 -688 -1597 688
rect -1563 -688 -1551 688
rect -1609 -700 -1551 -688
rect -1451 688 -1393 700
rect -1451 -688 -1439 688
rect -1405 -688 -1393 688
rect -1451 -700 -1393 -688
rect -1293 688 -1235 700
rect -1293 -688 -1281 688
rect -1247 -688 -1235 688
rect -1293 -700 -1235 -688
rect -1135 688 -1077 700
rect -1135 -688 -1123 688
rect -1089 -688 -1077 688
rect -1135 -700 -1077 -688
rect -977 688 -919 700
rect -977 -688 -965 688
rect -931 -688 -919 688
rect -977 -700 -919 -688
rect -819 688 -761 700
rect -819 -688 -807 688
rect -773 -688 -761 688
rect -819 -700 -761 -688
rect -661 688 -603 700
rect -661 -688 -649 688
rect -615 -688 -603 688
rect -661 -700 -603 -688
rect -503 688 -445 700
rect -503 -688 -491 688
rect -457 -688 -445 688
rect -503 -700 -445 -688
rect -345 688 -287 700
rect -345 -688 -333 688
rect -299 -688 -287 688
rect -345 -700 -287 -688
rect -187 688 -129 700
rect -187 -688 -175 688
rect -141 -688 -129 688
rect -187 -700 -129 -688
rect -29 688 29 700
rect -29 -688 -17 688
rect 17 -688 29 688
rect -29 -700 29 -688
rect 129 688 187 700
rect 129 -688 141 688
rect 175 -688 187 688
rect 129 -700 187 -688
rect 287 688 345 700
rect 287 -688 299 688
rect 333 -688 345 688
rect 287 -700 345 -688
rect 445 688 503 700
rect 445 -688 457 688
rect 491 -688 503 688
rect 445 -700 503 -688
rect 603 688 661 700
rect 603 -688 615 688
rect 649 -688 661 688
rect 603 -700 661 -688
rect 761 688 819 700
rect 761 -688 773 688
rect 807 -688 819 688
rect 761 -700 819 -688
rect 919 688 977 700
rect 919 -688 931 688
rect 965 -688 977 688
rect 919 -700 977 -688
rect 1077 688 1135 700
rect 1077 -688 1089 688
rect 1123 -688 1135 688
rect 1077 -700 1135 -688
rect 1235 688 1293 700
rect 1235 -688 1247 688
rect 1281 -688 1293 688
rect 1235 -700 1293 -688
rect 1393 688 1451 700
rect 1393 -688 1405 688
rect 1439 -688 1451 688
rect 1393 -700 1451 -688
rect 1551 688 1609 700
rect 1551 -688 1563 688
rect 1597 -688 1609 688
rect 1551 -700 1609 -688
rect 1709 688 1767 700
rect 1709 -688 1721 688
rect 1755 -688 1767 688
rect 1709 -700 1767 -688
rect 1867 688 1925 700
rect 1867 -688 1879 688
rect 1913 -688 1925 688
rect 1867 -700 1925 -688
rect 2025 688 2083 700
rect 2025 -688 2037 688
rect 2071 -688 2083 688
rect 2025 -700 2083 -688
rect 2183 688 2241 700
rect 2183 -688 2195 688
rect 2229 -688 2241 688
rect 2183 -700 2241 -688
rect 2341 688 2399 700
rect 2341 -688 2353 688
rect 2387 -688 2399 688
rect 2341 -700 2399 -688
rect 2499 688 2557 700
rect 2499 -688 2511 688
rect 2545 -688 2557 688
rect 2499 -700 2557 -688
rect 2657 688 2715 700
rect 2657 -688 2669 688
rect 2703 -688 2715 688
rect 2657 -700 2715 -688
rect 2815 688 2873 700
rect 2815 -688 2827 688
rect 2861 -688 2873 688
rect 2815 -700 2873 -688
rect 2973 688 3031 700
rect 2973 -688 2985 688
rect 3019 -688 3031 688
rect 2973 -700 3031 -688
rect 3131 688 3189 700
rect 3131 -688 3143 688
rect 3177 -688 3189 688
rect 3131 -700 3189 -688
rect 3289 688 3347 700
rect 3289 -688 3301 688
rect 3335 -688 3347 688
rect 3289 -700 3347 -688
rect 3447 688 3505 700
rect 3447 -688 3459 688
rect 3493 -688 3505 688
rect 3447 -700 3505 -688
rect 3605 688 3663 700
rect 3605 -688 3617 688
rect 3651 -688 3663 688
rect 3605 -700 3663 -688
rect 3763 688 3821 700
rect 3763 -688 3775 688
rect 3809 -688 3821 688
rect 3763 -700 3821 -688
rect 3921 688 3979 700
rect 3921 -688 3933 688
rect 3967 -688 3979 688
rect 3921 -700 3979 -688
rect 4079 688 4137 700
rect 4079 -688 4091 688
rect 4125 -688 4137 688
rect 4079 -700 4137 -688
rect 4237 688 4295 700
rect 4237 -688 4249 688
rect 4283 -688 4295 688
rect 4237 -700 4295 -688
rect 4395 688 4453 700
rect 4395 -688 4407 688
rect 4441 -688 4453 688
rect 4395 -700 4453 -688
rect 4553 688 4611 700
rect 4553 -688 4565 688
rect 4599 -688 4611 688
rect 4553 -700 4611 -688
rect 4711 688 4769 700
rect 4711 -688 4723 688
rect 4757 -688 4769 688
rect 4711 -700 4769 -688
rect 4869 688 4927 700
rect 4869 -688 4881 688
rect 4915 -688 4927 688
rect 4869 -700 4927 -688
rect 5027 688 5085 700
rect 5027 -688 5039 688
rect 5073 -688 5085 688
rect 5027 -700 5085 -688
rect 5185 688 5243 700
rect 5185 -688 5197 688
rect 5231 -688 5243 688
rect 5185 -700 5243 -688
rect 5343 688 5401 700
rect 5343 -688 5355 688
rect 5389 -688 5401 688
rect 5343 -700 5401 -688
rect 5501 688 5559 700
rect 5501 -688 5513 688
rect 5547 -688 5559 688
rect 5501 -700 5559 -688
rect 5659 688 5717 700
rect 5659 -688 5671 688
rect 5705 -688 5717 688
rect 5659 -700 5717 -688
rect 5817 688 5875 700
rect 5817 -688 5829 688
rect 5863 -688 5875 688
rect 5817 -700 5875 -688
rect 5975 688 6033 700
rect 5975 -688 5987 688
rect 6021 -688 6033 688
rect 5975 -700 6033 -688
rect 6133 688 6191 700
rect 6133 -688 6145 688
rect 6179 -688 6191 688
rect 6133 -700 6191 -688
rect 6291 688 6349 700
rect 6291 -688 6303 688
rect 6337 -688 6349 688
rect 6291 -700 6349 -688
rect 6449 688 6507 700
rect 6449 -688 6461 688
rect 6495 -688 6507 688
rect 6449 -700 6507 -688
rect 6607 688 6665 700
rect 6607 -688 6619 688
rect 6653 -688 6665 688
rect 6607 -700 6665 -688
rect 6765 688 6823 700
rect 6765 -688 6777 688
rect 6811 -688 6823 688
rect 6765 -700 6823 -688
rect 6923 688 6981 700
rect 6923 -688 6935 688
rect 6969 -688 6981 688
rect 6923 -700 6981 -688
<< mvndiffc >>
rect -6969 -688 -6935 688
rect -6811 -688 -6777 688
rect -6653 -688 -6619 688
rect -6495 -688 -6461 688
rect -6337 -688 -6303 688
rect -6179 -688 -6145 688
rect -6021 -688 -5987 688
rect -5863 -688 -5829 688
rect -5705 -688 -5671 688
rect -5547 -688 -5513 688
rect -5389 -688 -5355 688
rect -5231 -688 -5197 688
rect -5073 -688 -5039 688
rect -4915 -688 -4881 688
rect -4757 -688 -4723 688
rect -4599 -688 -4565 688
rect -4441 -688 -4407 688
rect -4283 -688 -4249 688
rect -4125 -688 -4091 688
rect -3967 -688 -3933 688
rect -3809 -688 -3775 688
rect -3651 -688 -3617 688
rect -3493 -688 -3459 688
rect -3335 -688 -3301 688
rect -3177 -688 -3143 688
rect -3019 -688 -2985 688
rect -2861 -688 -2827 688
rect -2703 -688 -2669 688
rect -2545 -688 -2511 688
rect -2387 -688 -2353 688
rect -2229 -688 -2195 688
rect -2071 -688 -2037 688
rect -1913 -688 -1879 688
rect -1755 -688 -1721 688
rect -1597 -688 -1563 688
rect -1439 -688 -1405 688
rect -1281 -688 -1247 688
rect -1123 -688 -1089 688
rect -965 -688 -931 688
rect -807 -688 -773 688
rect -649 -688 -615 688
rect -491 -688 -457 688
rect -333 -688 -299 688
rect -175 -688 -141 688
rect -17 -688 17 688
rect 141 -688 175 688
rect 299 -688 333 688
rect 457 -688 491 688
rect 615 -688 649 688
rect 773 -688 807 688
rect 931 -688 965 688
rect 1089 -688 1123 688
rect 1247 -688 1281 688
rect 1405 -688 1439 688
rect 1563 -688 1597 688
rect 1721 -688 1755 688
rect 1879 -688 1913 688
rect 2037 -688 2071 688
rect 2195 -688 2229 688
rect 2353 -688 2387 688
rect 2511 -688 2545 688
rect 2669 -688 2703 688
rect 2827 -688 2861 688
rect 2985 -688 3019 688
rect 3143 -688 3177 688
rect 3301 -688 3335 688
rect 3459 -688 3493 688
rect 3617 -688 3651 688
rect 3775 -688 3809 688
rect 3933 -688 3967 688
rect 4091 -688 4125 688
rect 4249 -688 4283 688
rect 4407 -688 4441 688
rect 4565 -688 4599 688
rect 4723 -688 4757 688
rect 4881 -688 4915 688
rect 5039 -688 5073 688
rect 5197 -688 5231 688
rect 5355 -688 5389 688
rect 5513 -688 5547 688
rect 5671 -688 5705 688
rect 5829 -688 5863 688
rect 5987 -688 6021 688
rect 6145 -688 6179 688
rect 6303 -688 6337 688
rect 6461 -688 6495 688
rect 6619 -688 6653 688
rect 6777 -688 6811 688
rect 6935 -688 6969 688
<< poly >>
rect -6923 772 -6823 788
rect -6923 738 -6907 772
rect -6839 738 -6823 772
rect -6923 700 -6823 738
rect -6765 772 -6665 788
rect -6765 738 -6749 772
rect -6681 738 -6665 772
rect -6765 700 -6665 738
rect -6607 772 -6507 788
rect -6607 738 -6591 772
rect -6523 738 -6507 772
rect -6607 700 -6507 738
rect -6449 772 -6349 788
rect -6449 738 -6433 772
rect -6365 738 -6349 772
rect -6449 700 -6349 738
rect -6291 772 -6191 788
rect -6291 738 -6275 772
rect -6207 738 -6191 772
rect -6291 700 -6191 738
rect -6133 772 -6033 788
rect -6133 738 -6117 772
rect -6049 738 -6033 772
rect -6133 700 -6033 738
rect -5975 772 -5875 788
rect -5975 738 -5959 772
rect -5891 738 -5875 772
rect -5975 700 -5875 738
rect -5817 772 -5717 788
rect -5817 738 -5801 772
rect -5733 738 -5717 772
rect -5817 700 -5717 738
rect -5659 772 -5559 788
rect -5659 738 -5643 772
rect -5575 738 -5559 772
rect -5659 700 -5559 738
rect -5501 772 -5401 788
rect -5501 738 -5485 772
rect -5417 738 -5401 772
rect -5501 700 -5401 738
rect -5343 772 -5243 788
rect -5343 738 -5327 772
rect -5259 738 -5243 772
rect -5343 700 -5243 738
rect -5185 772 -5085 788
rect -5185 738 -5169 772
rect -5101 738 -5085 772
rect -5185 700 -5085 738
rect -5027 772 -4927 788
rect -5027 738 -5011 772
rect -4943 738 -4927 772
rect -5027 700 -4927 738
rect -4869 772 -4769 788
rect -4869 738 -4853 772
rect -4785 738 -4769 772
rect -4869 700 -4769 738
rect -4711 772 -4611 788
rect -4711 738 -4695 772
rect -4627 738 -4611 772
rect -4711 700 -4611 738
rect -4553 772 -4453 788
rect -4553 738 -4537 772
rect -4469 738 -4453 772
rect -4553 700 -4453 738
rect -4395 772 -4295 788
rect -4395 738 -4379 772
rect -4311 738 -4295 772
rect -4395 700 -4295 738
rect -4237 772 -4137 788
rect -4237 738 -4221 772
rect -4153 738 -4137 772
rect -4237 700 -4137 738
rect -4079 772 -3979 788
rect -4079 738 -4063 772
rect -3995 738 -3979 772
rect -4079 700 -3979 738
rect -3921 772 -3821 788
rect -3921 738 -3905 772
rect -3837 738 -3821 772
rect -3921 700 -3821 738
rect -3763 772 -3663 788
rect -3763 738 -3747 772
rect -3679 738 -3663 772
rect -3763 700 -3663 738
rect -3605 772 -3505 788
rect -3605 738 -3589 772
rect -3521 738 -3505 772
rect -3605 700 -3505 738
rect -3447 772 -3347 788
rect -3447 738 -3431 772
rect -3363 738 -3347 772
rect -3447 700 -3347 738
rect -3289 772 -3189 788
rect -3289 738 -3273 772
rect -3205 738 -3189 772
rect -3289 700 -3189 738
rect -3131 772 -3031 788
rect -3131 738 -3115 772
rect -3047 738 -3031 772
rect -3131 700 -3031 738
rect -2973 772 -2873 788
rect -2973 738 -2957 772
rect -2889 738 -2873 772
rect -2973 700 -2873 738
rect -2815 772 -2715 788
rect -2815 738 -2799 772
rect -2731 738 -2715 772
rect -2815 700 -2715 738
rect -2657 772 -2557 788
rect -2657 738 -2641 772
rect -2573 738 -2557 772
rect -2657 700 -2557 738
rect -2499 772 -2399 788
rect -2499 738 -2483 772
rect -2415 738 -2399 772
rect -2499 700 -2399 738
rect -2341 772 -2241 788
rect -2341 738 -2325 772
rect -2257 738 -2241 772
rect -2341 700 -2241 738
rect -2183 772 -2083 788
rect -2183 738 -2167 772
rect -2099 738 -2083 772
rect -2183 700 -2083 738
rect -2025 772 -1925 788
rect -2025 738 -2009 772
rect -1941 738 -1925 772
rect -2025 700 -1925 738
rect -1867 772 -1767 788
rect -1867 738 -1851 772
rect -1783 738 -1767 772
rect -1867 700 -1767 738
rect -1709 772 -1609 788
rect -1709 738 -1693 772
rect -1625 738 -1609 772
rect -1709 700 -1609 738
rect -1551 772 -1451 788
rect -1551 738 -1535 772
rect -1467 738 -1451 772
rect -1551 700 -1451 738
rect -1393 772 -1293 788
rect -1393 738 -1377 772
rect -1309 738 -1293 772
rect -1393 700 -1293 738
rect -1235 772 -1135 788
rect -1235 738 -1219 772
rect -1151 738 -1135 772
rect -1235 700 -1135 738
rect -1077 772 -977 788
rect -1077 738 -1061 772
rect -993 738 -977 772
rect -1077 700 -977 738
rect -919 772 -819 788
rect -919 738 -903 772
rect -835 738 -819 772
rect -919 700 -819 738
rect -761 772 -661 788
rect -761 738 -745 772
rect -677 738 -661 772
rect -761 700 -661 738
rect -603 772 -503 788
rect -603 738 -587 772
rect -519 738 -503 772
rect -603 700 -503 738
rect -445 772 -345 788
rect -445 738 -429 772
rect -361 738 -345 772
rect -445 700 -345 738
rect -287 772 -187 788
rect -287 738 -271 772
rect -203 738 -187 772
rect -287 700 -187 738
rect -129 772 -29 788
rect -129 738 -113 772
rect -45 738 -29 772
rect -129 700 -29 738
rect 29 772 129 788
rect 29 738 45 772
rect 113 738 129 772
rect 29 700 129 738
rect 187 772 287 788
rect 187 738 203 772
rect 271 738 287 772
rect 187 700 287 738
rect 345 772 445 788
rect 345 738 361 772
rect 429 738 445 772
rect 345 700 445 738
rect 503 772 603 788
rect 503 738 519 772
rect 587 738 603 772
rect 503 700 603 738
rect 661 772 761 788
rect 661 738 677 772
rect 745 738 761 772
rect 661 700 761 738
rect 819 772 919 788
rect 819 738 835 772
rect 903 738 919 772
rect 819 700 919 738
rect 977 772 1077 788
rect 977 738 993 772
rect 1061 738 1077 772
rect 977 700 1077 738
rect 1135 772 1235 788
rect 1135 738 1151 772
rect 1219 738 1235 772
rect 1135 700 1235 738
rect 1293 772 1393 788
rect 1293 738 1309 772
rect 1377 738 1393 772
rect 1293 700 1393 738
rect 1451 772 1551 788
rect 1451 738 1467 772
rect 1535 738 1551 772
rect 1451 700 1551 738
rect 1609 772 1709 788
rect 1609 738 1625 772
rect 1693 738 1709 772
rect 1609 700 1709 738
rect 1767 772 1867 788
rect 1767 738 1783 772
rect 1851 738 1867 772
rect 1767 700 1867 738
rect 1925 772 2025 788
rect 1925 738 1941 772
rect 2009 738 2025 772
rect 1925 700 2025 738
rect 2083 772 2183 788
rect 2083 738 2099 772
rect 2167 738 2183 772
rect 2083 700 2183 738
rect 2241 772 2341 788
rect 2241 738 2257 772
rect 2325 738 2341 772
rect 2241 700 2341 738
rect 2399 772 2499 788
rect 2399 738 2415 772
rect 2483 738 2499 772
rect 2399 700 2499 738
rect 2557 772 2657 788
rect 2557 738 2573 772
rect 2641 738 2657 772
rect 2557 700 2657 738
rect 2715 772 2815 788
rect 2715 738 2731 772
rect 2799 738 2815 772
rect 2715 700 2815 738
rect 2873 772 2973 788
rect 2873 738 2889 772
rect 2957 738 2973 772
rect 2873 700 2973 738
rect 3031 772 3131 788
rect 3031 738 3047 772
rect 3115 738 3131 772
rect 3031 700 3131 738
rect 3189 772 3289 788
rect 3189 738 3205 772
rect 3273 738 3289 772
rect 3189 700 3289 738
rect 3347 772 3447 788
rect 3347 738 3363 772
rect 3431 738 3447 772
rect 3347 700 3447 738
rect 3505 772 3605 788
rect 3505 738 3521 772
rect 3589 738 3605 772
rect 3505 700 3605 738
rect 3663 772 3763 788
rect 3663 738 3679 772
rect 3747 738 3763 772
rect 3663 700 3763 738
rect 3821 772 3921 788
rect 3821 738 3837 772
rect 3905 738 3921 772
rect 3821 700 3921 738
rect 3979 772 4079 788
rect 3979 738 3995 772
rect 4063 738 4079 772
rect 3979 700 4079 738
rect 4137 772 4237 788
rect 4137 738 4153 772
rect 4221 738 4237 772
rect 4137 700 4237 738
rect 4295 772 4395 788
rect 4295 738 4311 772
rect 4379 738 4395 772
rect 4295 700 4395 738
rect 4453 772 4553 788
rect 4453 738 4469 772
rect 4537 738 4553 772
rect 4453 700 4553 738
rect 4611 772 4711 788
rect 4611 738 4627 772
rect 4695 738 4711 772
rect 4611 700 4711 738
rect 4769 772 4869 788
rect 4769 738 4785 772
rect 4853 738 4869 772
rect 4769 700 4869 738
rect 4927 772 5027 788
rect 4927 738 4943 772
rect 5011 738 5027 772
rect 4927 700 5027 738
rect 5085 772 5185 788
rect 5085 738 5101 772
rect 5169 738 5185 772
rect 5085 700 5185 738
rect 5243 772 5343 788
rect 5243 738 5259 772
rect 5327 738 5343 772
rect 5243 700 5343 738
rect 5401 772 5501 788
rect 5401 738 5417 772
rect 5485 738 5501 772
rect 5401 700 5501 738
rect 5559 772 5659 788
rect 5559 738 5575 772
rect 5643 738 5659 772
rect 5559 700 5659 738
rect 5717 772 5817 788
rect 5717 738 5733 772
rect 5801 738 5817 772
rect 5717 700 5817 738
rect 5875 772 5975 788
rect 5875 738 5891 772
rect 5959 738 5975 772
rect 5875 700 5975 738
rect 6033 772 6133 788
rect 6033 738 6049 772
rect 6117 738 6133 772
rect 6033 700 6133 738
rect 6191 772 6291 788
rect 6191 738 6207 772
rect 6275 738 6291 772
rect 6191 700 6291 738
rect 6349 772 6449 788
rect 6349 738 6365 772
rect 6433 738 6449 772
rect 6349 700 6449 738
rect 6507 772 6607 788
rect 6507 738 6523 772
rect 6591 738 6607 772
rect 6507 700 6607 738
rect 6665 772 6765 788
rect 6665 738 6681 772
rect 6749 738 6765 772
rect 6665 700 6765 738
rect 6823 772 6923 788
rect 6823 738 6839 772
rect 6907 738 6923 772
rect 6823 700 6923 738
rect -6923 -738 -6823 -700
rect -6923 -772 -6907 -738
rect -6839 -772 -6823 -738
rect -6923 -788 -6823 -772
rect -6765 -738 -6665 -700
rect -6765 -772 -6749 -738
rect -6681 -772 -6665 -738
rect -6765 -788 -6665 -772
rect -6607 -738 -6507 -700
rect -6607 -772 -6591 -738
rect -6523 -772 -6507 -738
rect -6607 -788 -6507 -772
rect -6449 -738 -6349 -700
rect -6449 -772 -6433 -738
rect -6365 -772 -6349 -738
rect -6449 -788 -6349 -772
rect -6291 -738 -6191 -700
rect -6291 -772 -6275 -738
rect -6207 -772 -6191 -738
rect -6291 -788 -6191 -772
rect -6133 -738 -6033 -700
rect -6133 -772 -6117 -738
rect -6049 -772 -6033 -738
rect -6133 -788 -6033 -772
rect -5975 -738 -5875 -700
rect -5975 -772 -5959 -738
rect -5891 -772 -5875 -738
rect -5975 -788 -5875 -772
rect -5817 -738 -5717 -700
rect -5817 -772 -5801 -738
rect -5733 -772 -5717 -738
rect -5817 -788 -5717 -772
rect -5659 -738 -5559 -700
rect -5659 -772 -5643 -738
rect -5575 -772 -5559 -738
rect -5659 -788 -5559 -772
rect -5501 -738 -5401 -700
rect -5501 -772 -5485 -738
rect -5417 -772 -5401 -738
rect -5501 -788 -5401 -772
rect -5343 -738 -5243 -700
rect -5343 -772 -5327 -738
rect -5259 -772 -5243 -738
rect -5343 -788 -5243 -772
rect -5185 -738 -5085 -700
rect -5185 -772 -5169 -738
rect -5101 -772 -5085 -738
rect -5185 -788 -5085 -772
rect -5027 -738 -4927 -700
rect -5027 -772 -5011 -738
rect -4943 -772 -4927 -738
rect -5027 -788 -4927 -772
rect -4869 -738 -4769 -700
rect -4869 -772 -4853 -738
rect -4785 -772 -4769 -738
rect -4869 -788 -4769 -772
rect -4711 -738 -4611 -700
rect -4711 -772 -4695 -738
rect -4627 -772 -4611 -738
rect -4711 -788 -4611 -772
rect -4553 -738 -4453 -700
rect -4553 -772 -4537 -738
rect -4469 -772 -4453 -738
rect -4553 -788 -4453 -772
rect -4395 -738 -4295 -700
rect -4395 -772 -4379 -738
rect -4311 -772 -4295 -738
rect -4395 -788 -4295 -772
rect -4237 -738 -4137 -700
rect -4237 -772 -4221 -738
rect -4153 -772 -4137 -738
rect -4237 -788 -4137 -772
rect -4079 -738 -3979 -700
rect -4079 -772 -4063 -738
rect -3995 -772 -3979 -738
rect -4079 -788 -3979 -772
rect -3921 -738 -3821 -700
rect -3921 -772 -3905 -738
rect -3837 -772 -3821 -738
rect -3921 -788 -3821 -772
rect -3763 -738 -3663 -700
rect -3763 -772 -3747 -738
rect -3679 -772 -3663 -738
rect -3763 -788 -3663 -772
rect -3605 -738 -3505 -700
rect -3605 -772 -3589 -738
rect -3521 -772 -3505 -738
rect -3605 -788 -3505 -772
rect -3447 -738 -3347 -700
rect -3447 -772 -3431 -738
rect -3363 -772 -3347 -738
rect -3447 -788 -3347 -772
rect -3289 -738 -3189 -700
rect -3289 -772 -3273 -738
rect -3205 -772 -3189 -738
rect -3289 -788 -3189 -772
rect -3131 -738 -3031 -700
rect -3131 -772 -3115 -738
rect -3047 -772 -3031 -738
rect -3131 -788 -3031 -772
rect -2973 -738 -2873 -700
rect -2973 -772 -2957 -738
rect -2889 -772 -2873 -738
rect -2973 -788 -2873 -772
rect -2815 -738 -2715 -700
rect -2815 -772 -2799 -738
rect -2731 -772 -2715 -738
rect -2815 -788 -2715 -772
rect -2657 -738 -2557 -700
rect -2657 -772 -2641 -738
rect -2573 -772 -2557 -738
rect -2657 -788 -2557 -772
rect -2499 -738 -2399 -700
rect -2499 -772 -2483 -738
rect -2415 -772 -2399 -738
rect -2499 -788 -2399 -772
rect -2341 -738 -2241 -700
rect -2341 -772 -2325 -738
rect -2257 -772 -2241 -738
rect -2341 -788 -2241 -772
rect -2183 -738 -2083 -700
rect -2183 -772 -2167 -738
rect -2099 -772 -2083 -738
rect -2183 -788 -2083 -772
rect -2025 -738 -1925 -700
rect -2025 -772 -2009 -738
rect -1941 -772 -1925 -738
rect -2025 -788 -1925 -772
rect -1867 -738 -1767 -700
rect -1867 -772 -1851 -738
rect -1783 -772 -1767 -738
rect -1867 -788 -1767 -772
rect -1709 -738 -1609 -700
rect -1709 -772 -1693 -738
rect -1625 -772 -1609 -738
rect -1709 -788 -1609 -772
rect -1551 -738 -1451 -700
rect -1551 -772 -1535 -738
rect -1467 -772 -1451 -738
rect -1551 -788 -1451 -772
rect -1393 -738 -1293 -700
rect -1393 -772 -1377 -738
rect -1309 -772 -1293 -738
rect -1393 -788 -1293 -772
rect -1235 -738 -1135 -700
rect -1235 -772 -1219 -738
rect -1151 -772 -1135 -738
rect -1235 -788 -1135 -772
rect -1077 -738 -977 -700
rect -1077 -772 -1061 -738
rect -993 -772 -977 -738
rect -1077 -788 -977 -772
rect -919 -738 -819 -700
rect -919 -772 -903 -738
rect -835 -772 -819 -738
rect -919 -788 -819 -772
rect -761 -738 -661 -700
rect -761 -772 -745 -738
rect -677 -772 -661 -738
rect -761 -788 -661 -772
rect -603 -738 -503 -700
rect -603 -772 -587 -738
rect -519 -772 -503 -738
rect -603 -788 -503 -772
rect -445 -738 -345 -700
rect -445 -772 -429 -738
rect -361 -772 -345 -738
rect -445 -788 -345 -772
rect -287 -738 -187 -700
rect -287 -772 -271 -738
rect -203 -772 -187 -738
rect -287 -788 -187 -772
rect -129 -738 -29 -700
rect -129 -772 -113 -738
rect -45 -772 -29 -738
rect -129 -788 -29 -772
rect 29 -738 129 -700
rect 29 -772 45 -738
rect 113 -772 129 -738
rect 29 -788 129 -772
rect 187 -738 287 -700
rect 187 -772 203 -738
rect 271 -772 287 -738
rect 187 -788 287 -772
rect 345 -738 445 -700
rect 345 -772 361 -738
rect 429 -772 445 -738
rect 345 -788 445 -772
rect 503 -738 603 -700
rect 503 -772 519 -738
rect 587 -772 603 -738
rect 503 -788 603 -772
rect 661 -738 761 -700
rect 661 -772 677 -738
rect 745 -772 761 -738
rect 661 -788 761 -772
rect 819 -738 919 -700
rect 819 -772 835 -738
rect 903 -772 919 -738
rect 819 -788 919 -772
rect 977 -738 1077 -700
rect 977 -772 993 -738
rect 1061 -772 1077 -738
rect 977 -788 1077 -772
rect 1135 -738 1235 -700
rect 1135 -772 1151 -738
rect 1219 -772 1235 -738
rect 1135 -788 1235 -772
rect 1293 -738 1393 -700
rect 1293 -772 1309 -738
rect 1377 -772 1393 -738
rect 1293 -788 1393 -772
rect 1451 -738 1551 -700
rect 1451 -772 1467 -738
rect 1535 -772 1551 -738
rect 1451 -788 1551 -772
rect 1609 -738 1709 -700
rect 1609 -772 1625 -738
rect 1693 -772 1709 -738
rect 1609 -788 1709 -772
rect 1767 -738 1867 -700
rect 1767 -772 1783 -738
rect 1851 -772 1867 -738
rect 1767 -788 1867 -772
rect 1925 -738 2025 -700
rect 1925 -772 1941 -738
rect 2009 -772 2025 -738
rect 1925 -788 2025 -772
rect 2083 -738 2183 -700
rect 2083 -772 2099 -738
rect 2167 -772 2183 -738
rect 2083 -788 2183 -772
rect 2241 -738 2341 -700
rect 2241 -772 2257 -738
rect 2325 -772 2341 -738
rect 2241 -788 2341 -772
rect 2399 -738 2499 -700
rect 2399 -772 2415 -738
rect 2483 -772 2499 -738
rect 2399 -788 2499 -772
rect 2557 -738 2657 -700
rect 2557 -772 2573 -738
rect 2641 -772 2657 -738
rect 2557 -788 2657 -772
rect 2715 -738 2815 -700
rect 2715 -772 2731 -738
rect 2799 -772 2815 -738
rect 2715 -788 2815 -772
rect 2873 -738 2973 -700
rect 2873 -772 2889 -738
rect 2957 -772 2973 -738
rect 2873 -788 2973 -772
rect 3031 -738 3131 -700
rect 3031 -772 3047 -738
rect 3115 -772 3131 -738
rect 3031 -788 3131 -772
rect 3189 -738 3289 -700
rect 3189 -772 3205 -738
rect 3273 -772 3289 -738
rect 3189 -788 3289 -772
rect 3347 -738 3447 -700
rect 3347 -772 3363 -738
rect 3431 -772 3447 -738
rect 3347 -788 3447 -772
rect 3505 -738 3605 -700
rect 3505 -772 3521 -738
rect 3589 -772 3605 -738
rect 3505 -788 3605 -772
rect 3663 -738 3763 -700
rect 3663 -772 3679 -738
rect 3747 -772 3763 -738
rect 3663 -788 3763 -772
rect 3821 -738 3921 -700
rect 3821 -772 3837 -738
rect 3905 -772 3921 -738
rect 3821 -788 3921 -772
rect 3979 -738 4079 -700
rect 3979 -772 3995 -738
rect 4063 -772 4079 -738
rect 3979 -788 4079 -772
rect 4137 -738 4237 -700
rect 4137 -772 4153 -738
rect 4221 -772 4237 -738
rect 4137 -788 4237 -772
rect 4295 -738 4395 -700
rect 4295 -772 4311 -738
rect 4379 -772 4395 -738
rect 4295 -788 4395 -772
rect 4453 -738 4553 -700
rect 4453 -772 4469 -738
rect 4537 -772 4553 -738
rect 4453 -788 4553 -772
rect 4611 -738 4711 -700
rect 4611 -772 4627 -738
rect 4695 -772 4711 -738
rect 4611 -788 4711 -772
rect 4769 -738 4869 -700
rect 4769 -772 4785 -738
rect 4853 -772 4869 -738
rect 4769 -788 4869 -772
rect 4927 -738 5027 -700
rect 4927 -772 4943 -738
rect 5011 -772 5027 -738
rect 4927 -788 5027 -772
rect 5085 -738 5185 -700
rect 5085 -772 5101 -738
rect 5169 -772 5185 -738
rect 5085 -788 5185 -772
rect 5243 -738 5343 -700
rect 5243 -772 5259 -738
rect 5327 -772 5343 -738
rect 5243 -788 5343 -772
rect 5401 -738 5501 -700
rect 5401 -772 5417 -738
rect 5485 -772 5501 -738
rect 5401 -788 5501 -772
rect 5559 -738 5659 -700
rect 5559 -772 5575 -738
rect 5643 -772 5659 -738
rect 5559 -788 5659 -772
rect 5717 -738 5817 -700
rect 5717 -772 5733 -738
rect 5801 -772 5817 -738
rect 5717 -788 5817 -772
rect 5875 -738 5975 -700
rect 5875 -772 5891 -738
rect 5959 -772 5975 -738
rect 5875 -788 5975 -772
rect 6033 -738 6133 -700
rect 6033 -772 6049 -738
rect 6117 -772 6133 -738
rect 6033 -788 6133 -772
rect 6191 -738 6291 -700
rect 6191 -772 6207 -738
rect 6275 -772 6291 -738
rect 6191 -788 6291 -772
rect 6349 -738 6449 -700
rect 6349 -772 6365 -738
rect 6433 -772 6449 -738
rect 6349 -788 6449 -772
rect 6507 -738 6607 -700
rect 6507 -772 6523 -738
rect 6591 -772 6607 -738
rect 6507 -788 6607 -772
rect 6665 -738 6765 -700
rect 6665 -772 6681 -738
rect 6749 -772 6765 -738
rect 6665 -788 6765 -772
rect 6823 -738 6923 -700
rect 6823 -772 6839 -738
rect 6907 -772 6923 -738
rect 6823 -788 6923 -772
<< polycont >>
rect -6907 738 -6839 772
rect -6749 738 -6681 772
rect -6591 738 -6523 772
rect -6433 738 -6365 772
rect -6275 738 -6207 772
rect -6117 738 -6049 772
rect -5959 738 -5891 772
rect -5801 738 -5733 772
rect -5643 738 -5575 772
rect -5485 738 -5417 772
rect -5327 738 -5259 772
rect -5169 738 -5101 772
rect -5011 738 -4943 772
rect -4853 738 -4785 772
rect -4695 738 -4627 772
rect -4537 738 -4469 772
rect -4379 738 -4311 772
rect -4221 738 -4153 772
rect -4063 738 -3995 772
rect -3905 738 -3837 772
rect -3747 738 -3679 772
rect -3589 738 -3521 772
rect -3431 738 -3363 772
rect -3273 738 -3205 772
rect -3115 738 -3047 772
rect -2957 738 -2889 772
rect -2799 738 -2731 772
rect -2641 738 -2573 772
rect -2483 738 -2415 772
rect -2325 738 -2257 772
rect -2167 738 -2099 772
rect -2009 738 -1941 772
rect -1851 738 -1783 772
rect -1693 738 -1625 772
rect -1535 738 -1467 772
rect -1377 738 -1309 772
rect -1219 738 -1151 772
rect -1061 738 -993 772
rect -903 738 -835 772
rect -745 738 -677 772
rect -587 738 -519 772
rect -429 738 -361 772
rect -271 738 -203 772
rect -113 738 -45 772
rect 45 738 113 772
rect 203 738 271 772
rect 361 738 429 772
rect 519 738 587 772
rect 677 738 745 772
rect 835 738 903 772
rect 993 738 1061 772
rect 1151 738 1219 772
rect 1309 738 1377 772
rect 1467 738 1535 772
rect 1625 738 1693 772
rect 1783 738 1851 772
rect 1941 738 2009 772
rect 2099 738 2167 772
rect 2257 738 2325 772
rect 2415 738 2483 772
rect 2573 738 2641 772
rect 2731 738 2799 772
rect 2889 738 2957 772
rect 3047 738 3115 772
rect 3205 738 3273 772
rect 3363 738 3431 772
rect 3521 738 3589 772
rect 3679 738 3747 772
rect 3837 738 3905 772
rect 3995 738 4063 772
rect 4153 738 4221 772
rect 4311 738 4379 772
rect 4469 738 4537 772
rect 4627 738 4695 772
rect 4785 738 4853 772
rect 4943 738 5011 772
rect 5101 738 5169 772
rect 5259 738 5327 772
rect 5417 738 5485 772
rect 5575 738 5643 772
rect 5733 738 5801 772
rect 5891 738 5959 772
rect 6049 738 6117 772
rect 6207 738 6275 772
rect 6365 738 6433 772
rect 6523 738 6591 772
rect 6681 738 6749 772
rect 6839 738 6907 772
rect -6907 -772 -6839 -738
rect -6749 -772 -6681 -738
rect -6591 -772 -6523 -738
rect -6433 -772 -6365 -738
rect -6275 -772 -6207 -738
rect -6117 -772 -6049 -738
rect -5959 -772 -5891 -738
rect -5801 -772 -5733 -738
rect -5643 -772 -5575 -738
rect -5485 -772 -5417 -738
rect -5327 -772 -5259 -738
rect -5169 -772 -5101 -738
rect -5011 -772 -4943 -738
rect -4853 -772 -4785 -738
rect -4695 -772 -4627 -738
rect -4537 -772 -4469 -738
rect -4379 -772 -4311 -738
rect -4221 -772 -4153 -738
rect -4063 -772 -3995 -738
rect -3905 -772 -3837 -738
rect -3747 -772 -3679 -738
rect -3589 -772 -3521 -738
rect -3431 -772 -3363 -738
rect -3273 -772 -3205 -738
rect -3115 -772 -3047 -738
rect -2957 -772 -2889 -738
rect -2799 -772 -2731 -738
rect -2641 -772 -2573 -738
rect -2483 -772 -2415 -738
rect -2325 -772 -2257 -738
rect -2167 -772 -2099 -738
rect -2009 -772 -1941 -738
rect -1851 -772 -1783 -738
rect -1693 -772 -1625 -738
rect -1535 -772 -1467 -738
rect -1377 -772 -1309 -738
rect -1219 -772 -1151 -738
rect -1061 -772 -993 -738
rect -903 -772 -835 -738
rect -745 -772 -677 -738
rect -587 -772 -519 -738
rect -429 -772 -361 -738
rect -271 -772 -203 -738
rect -113 -772 -45 -738
rect 45 -772 113 -738
rect 203 -772 271 -738
rect 361 -772 429 -738
rect 519 -772 587 -738
rect 677 -772 745 -738
rect 835 -772 903 -738
rect 993 -772 1061 -738
rect 1151 -772 1219 -738
rect 1309 -772 1377 -738
rect 1467 -772 1535 -738
rect 1625 -772 1693 -738
rect 1783 -772 1851 -738
rect 1941 -772 2009 -738
rect 2099 -772 2167 -738
rect 2257 -772 2325 -738
rect 2415 -772 2483 -738
rect 2573 -772 2641 -738
rect 2731 -772 2799 -738
rect 2889 -772 2957 -738
rect 3047 -772 3115 -738
rect 3205 -772 3273 -738
rect 3363 -772 3431 -738
rect 3521 -772 3589 -738
rect 3679 -772 3747 -738
rect 3837 -772 3905 -738
rect 3995 -772 4063 -738
rect 4153 -772 4221 -738
rect 4311 -772 4379 -738
rect 4469 -772 4537 -738
rect 4627 -772 4695 -738
rect 4785 -772 4853 -738
rect 4943 -772 5011 -738
rect 5101 -772 5169 -738
rect 5259 -772 5327 -738
rect 5417 -772 5485 -738
rect 5575 -772 5643 -738
rect 5733 -772 5801 -738
rect 5891 -772 5959 -738
rect 6049 -772 6117 -738
rect 6207 -772 6275 -738
rect 6365 -772 6433 -738
rect 6523 -772 6591 -738
rect 6681 -772 6749 -738
rect 6839 -772 6907 -738
<< locali >>
rect -6923 738 -6907 772
rect -6839 738 -6823 772
rect -6765 738 -6749 772
rect -6681 738 -6665 772
rect -6607 738 -6591 772
rect -6523 738 -6507 772
rect -6449 738 -6433 772
rect -6365 738 -6349 772
rect -6291 738 -6275 772
rect -6207 738 -6191 772
rect -6133 738 -6117 772
rect -6049 738 -6033 772
rect -5975 738 -5959 772
rect -5891 738 -5875 772
rect -5817 738 -5801 772
rect -5733 738 -5717 772
rect -5659 738 -5643 772
rect -5575 738 -5559 772
rect -5501 738 -5485 772
rect -5417 738 -5401 772
rect -5343 738 -5327 772
rect -5259 738 -5243 772
rect -5185 738 -5169 772
rect -5101 738 -5085 772
rect -5027 738 -5011 772
rect -4943 738 -4927 772
rect -4869 738 -4853 772
rect -4785 738 -4769 772
rect -4711 738 -4695 772
rect -4627 738 -4611 772
rect -4553 738 -4537 772
rect -4469 738 -4453 772
rect -4395 738 -4379 772
rect -4311 738 -4295 772
rect -4237 738 -4221 772
rect -4153 738 -4137 772
rect -4079 738 -4063 772
rect -3995 738 -3979 772
rect -3921 738 -3905 772
rect -3837 738 -3821 772
rect -3763 738 -3747 772
rect -3679 738 -3663 772
rect -3605 738 -3589 772
rect -3521 738 -3505 772
rect -3447 738 -3431 772
rect -3363 738 -3347 772
rect -3289 738 -3273 772
rect -3205 738 -3189 772
rect -3131 738 -3115 772
rect -3047 738 -3031 772
rect -2973 738 -2957 772
rect -2889 738 -2873 772
rect -2815 738 -2799 772
rect -2731 738 -2715 772
rect -2657 738 -2641 772
rect -2573 738 -2557 772
rect -2499 738 -2483 772
rect -2415 738 -2399 772
rect -2341 738 -2325 772
rect -2257 738 -2241 772
rect -2183 738 -2167 772
rect -2099 738 -2083 772
rect -2025 738 -2009 772
rect -1941 738 -1925 772
rect -1867 738 -1851 772
rect -1783 738 -1767 772
rect -1709 738 -1693 772
rect -1625 738 -1609 772
rect -1551 738 -1535 772
rect -1467 738 -1451 772
rect -1393 738 -1377 772
rect -1309 738 -1293 772
rect -1235 738 -1219 772
rect -1151 738 -1135 772
rect -1077 738 -1061 772
rect -993 738 -977 772
rect -919 738 -903 772
rect -835 738 -819 772
rect -761 738 -745 772
rect -677 738 -661 772
rect -603 738 -587 772
rect -519 738 -503 772
rect -445 738 -429 772
rect -361 738 -345 772
rect -287 738 -271 772
rect -203 738 -187 772
rect -129 738 -113 772
rect -45 738 -29 772
rect 29 738 45 772
rect 113 738 129 772
rect 187 738 203 772
rect 271 738 287 772
rect 345 738 361 772
rect 429 738 445 772
rect 503 738 519 772
rect 587 738 603 772
rect 661 738 677 772
rect 745 738 761 772
rect 819 738 835 772
rect 903 738 919 772
rect 977 738 993 772
rect 1061 738 1077 772
rect 1135 738 1151 772
rect 1219 738 1235 772
rect 1293 738 1309 772
rect 1377 738 1393 772
rect 1451 738 1467 772
rect 1535 738 1551 772
rect 1609 738 1625 772
rect 1693 738 1709 772
rect 1767 738 1783 772
rect 1851 738 1867 772
rect 1925 738 1941 772
rect 2009 738 2025 772
rect 2083 738 2099 772
rect 2167 738 2183 772
rect 2241 738 2257 772
rect 2325 738 2341 772
rect 2399 738 2415 772
rect 2483 738 2499 772
rect 2557 738 2573 772
rect 2641 738 2657 772
rect 2715 738 2731 772
rect 2799 738 2815 772
rect 2873 738 2889 772
rect 2957 738 2973 772
rect 3031 738 3047 772
rect 3115 738 3131 772
rect 3189 738 3205 772
rect 3273 738 3289 772
rect 3347 738 3363 772
rect 3431 738 3447 772
rect 3505 738 3521 772
rect 3589 738 3605 772
rect 3663 738 3679 772
rect 3747 738 3763 772
rect 3821 738 3837 772
rect 3905 738 3921 772
rect 3979 738 3995 772
rect 4063 738 4079 772
rect 4137 738 4153 772
rect 4221 738 4237 772
rect 4295 738 4311 772
rect 4379 738 4395 772
rect 4453 738 4469 772
rect 4537 738 4553 772
rect 4611 738 4627 772
rect 4695 738 4711 772
rect 4769 738 4785 772
rect 4853 738 4869 772
rect 4927 738 4943 772
rect 5011 738 5027 772
rect 5085 738 5101 772
rect 5169 738 5185 772
rect 5243 738 5259 772
rect 5327 738 5343 772
rect 5401 738 5417 772
rect 5485 738 5501 772
rect 5559 738 5575 772
rect 5643 738 5659 772
rect 5717 738 5733 772
rect 5801 738 5817 772
rect 5875 738 5891 772
rect 5959 738 5975 772
rect 6033 738 6049 772
rect 6117 738 6133 772
rect 6191 738 6207 772
rect 6275 738 6291 772
rect 6349 738 6365 772
rect 6433 738 6449 772
rect 6507 738 6523 772
rect 6591 738 6607 772
rect 6665 738 6681 772
rect 6749 738 6765 772
rect 6823 738 6839 772
rect 6907 738 6923 772
rect -6969 688 -6935 704
rect -6969 -704 -6935 -688
rect -6811 688 -6777 704
rect -6811 -704 -6777 -688
rect -6653 688 -6619 704
rect -6653 -704 -6619 -688
rect -6495 688 -6461 704
rect -6495 -704 -6461 -688
rect -6337 688 -6303 704
rect -6337 -704 -6303 -688
rect -6179 688 -6145 704
rect -6179 -704 -6145 -688
rect -6021 688 -5987 704
rect -6021 -704 -5987 -688
rect -5863 688 -5829 704
rect -5863 -704 -5829 -688
rect -5705 688 -5671 704
rect -5705 -704 -5671 -688
rect -5547 688 -5513 704
rect -5547 -704 -5513 -688
rect -5389 688 -5355 704
rect -5389 -704 -5355 -688
rect -5231 688 -5197 704
rect -5231 -704 -5197 -688
rect -5073 688 -5039 704
rect -5073 -704 -5039 -688
rect -4915 688 -4881 704
rect -4915 -704 -4881 -688
rect -4757 688 -4723 704
rect -4757 -704 -4723 -688
rect -4599 688 -4565 704
rect -4599 -704 -4565 -688
rect -4441 688 -4407 704
rect -4441 -704 -4407 -688
rect -4283 688 -4249 704
rect -4283 -704 -4249 -688
rect -4125 688 -4091 704
rect -4125 -704 -4091 -688
rect -3967 688 -3933 704
rect -3967 -704 -3933 -688
rect -3809 688 -3775 704
rect -3809 -704 -3775 -688
rect -3651 688 -3617 704
rect -3651 -704 -3617 -688
rect -3493 688 -3459 704
rect -3493 -704 -3459 -688
rect -3335 688 -3301 704
rect -3335 -704 -3301 -688
rect -3177 688 -3143 704
rect -3177 -704 -3143 -688
rect -3019 688 -2985 704
rect -3019 -704 -2985 -688
rect -2861 688 -2827 704
rect -2861 -704 -2827 -688
rect -2703 688 -2669 704
rect -2703 -704 -2669 -688
rect -2545 688 -2511 704
rect -2545 -704 -2511 -688
rect -2387 688 -2353 704
rect -2387 -704 -2353 -688
rect -2229 688 -2195 704
rect -2229 -704 -2195 -688
rect -2071 688 -2037 704
rect -2071 -704 -2037 -688
rect -1913 688 -1879 704
rect -1913 -704 -1879 -688
rect -1755 688 -1721 704
rect -1755 -704 -1721 -688
rect -1597 688 -1563 704
rect -1597 -704 -1563 -688
rect -1439 688 -1405 704
rect -1439 -704 -1405 -688
rect -1281 688 -1247 704
rect -1281 -704 -1247 -688
rect -1123 688 -1089 704
rect -1123 -704 -1089 -688
rect -965 688 -931 704
rect -965 -704 -931 -688
rect -807 688 -773 704
rect -807 -704 -773 -688
rect -649 688 -615 704
rect -649 -704 -615 -688
rect -491 688 -457 704
rect -491 -704 -457 -688
rect -333 688 -299 704
rect -333 -704 -299 -688
rect -175 688 -141 704
rect -175 -704 -141 -688
rect -17 688 17 704
rect -17 -704 17 -688
rect 141 688 175 704
rect 141 -704 175 -688
rect 299 688 333 704
rect 299 -704 333 -688
rect 457 688 491 704
rect 457 -704 491 -688
rect 615 688 649 704
rect 615 -704 649 -688
rect 773 688 807 704
rect 773 -704 807 -688
rect 931 688 965 704
rect 931 -704 965 -688
rect 1089 688 1123 704
rect 1089 -704 1123 -688
rect 1247 688 1281 704
rect 1247 -704 1281 -688
rect 1405 688 1439 704
rect 1405 -704 1439 -688
rect 1563 688 1597 704
rect 1563 -704 1597 -688
rect 1721 688 1755 704
rect 1721 -704 1755 -688
rect 1879 688 1913 704
rect 1879 -704 1913 -688
rect 2037 688 2071 704
rect 2037 -704 2071 -688
rect 2195 688 2229 704
rect 2195 -704 2229 -688
rect 2353 688 2387 704
rect 2353 -704 2387 -688
rect 2511 688 2545 704
rect 2511 -704 2545 -688
rect 2669 688 2703 704
rect 2669 -704 2703 -688
rect 2827 688 2861 704
rect 2827 -704 2861 -688
rect 2985 688 3019 704
rect 2985 -704 3019 -688
rect 3143 688 3177 704
rect 3143 -704 3177 -688
rect 3301 688 3335 704
rect 3301 -704 3335 -688
rect 3459 688 3493 704
rect 3459 -704 3493 -688
rect 3617 688 3651 704
rect 3617 -704 3651 -688
rect 3775 688 3809 704
rect 3775 -704 3809 -688
rect 3933 688 3967 704
rect 3933 -704 3967 -688
rect 4091 688 4125 704
rect 4091 -704 4125 -688
rect 4249 688 4283 704
rect 4249 -704 4283 -688
rect 4407 688 4441 704
rect 4407 -704 4441 -688
rect 4565 688 4599 704
rect 4565 -704 4599 -688
rect 4723 688 4757 704
rect 4723 -704 4757 -688
rect 4881 688 4915 704
rect 4881 -704 4915 -688
rect 5039 688 5073 704
rect 5039 -704 5073 -688
rect 5197 688 5231 704
rect 5197 -704 5231 -688
rect 5355 688 5389 704
rect 5355 -704 5389 -688
rect 5513 688 5547 704
rect 5513 -704 5547 -688
rect 5671 688 5705 704
rect 5671 -704 5705 -688
rect 5829 688 5863 704
rect 5829 -704 5863 -688
rect 5987 688 6021 704
rect 5987 -704 6021 -688
rect 6145 688 6179 704
rect 6145 -704 6179 -688
rect 6303 688 6337 704
rect 6303 -704 6337 -688
rect 6461 688 6495 704
rect 6461 -704 6495 -688
rect 6619 688 6653 704
rect 6619 -704 6653 -688
rect 6777 688 6811 704
rect 6777 -704 6811 -688
rect 6935 688 6969 704
rect 6935 -704 6969 -688
rect -6923 -772 -6907 -738
rect -6839 -772 -6823 -738
rect -6765 -772 -6749 -738
rect -6681 -772 -6665 -738
rect -6607 -772 -6591 -738
rect -6523 -772 -6507 -738
rect -6449 -772 -6433 -738
rect -6365 -772 -6349 -738
rect -6291 -772 -6275 -738
rect -6207 -772 -6191 -738
rect -6133 -772 -6117 -738
rect -6049 -772 -6033 -738
rect -5975 -772 -5959 -738
rect -5891 -772 -5875 -738
rect -5817 -772 -5801 -738
rect -5733 -772 -5717 -738
rect -5659 -772 -5643 -738
rect -5575 -772 -5559 -738
rect -5501 -772 -5485 -738
rect -5417 -772 -5401 -738
rect -5343 -772 -5327 -738
rect -5259 -772 -5243 -738
rect -5185 -772 -5169 -738
rect -5101 -772 -5085 -738
rect -5027 -772 -5011 -738
rect -4943 -772 -4927 -738
rect -4869 -772 -4853 -738
rect -4785 -772 -4769 -738
rect -4711 -772 -4695 -738
rect -4627 -772 -4611 -738
rect -4553 -772 -4537 -738
rect -4469 -772 -4453 -738
rect -4395 -772 -4379 -738
rect -4311 -772 -4295 -738
rect -4237 -772 -4221 -738
rect -4153 -772 -4137 -738
rect -4079 -772 -4063 -738
rect -3995 -772 -3979 -738
rect -3921 -772 -3905 -738
rect -3837 -772 -3821 -738
rect -3763 -772 -3747 -738
rect -3679 -772 -3663 -738
rect -3605 -772 -3589 -738
rect -3521 -772 -3505 -738
rect -3447 -772 -3431 -738
rect -3363 -772 -3347 -738
rect -3289 -772 -3273 -738
rect -3205 -772 -3189 -738
rect -3131 -772 -3115 -738
rect -3047 -772 -3031 -738
rect -2973 -772 -2957 -738
rect -2889 -772 -2873 -738
rect -2815 -772 -2799 -738
rect -2731 -772 -2715 -738
rect -2657 -772 -2641 -738
rect -2573 -772 -2557 -738
rect -2499 -772 -2483 -738
rect -2415 -772 -2399 -738
rect -2341 -772 -2325 -738
rect -2257 -772 -2241 -738
rect -2183 -772 -2167 -738
rect -2099 -772 -2083 -738
rect -2025 -772 -2009 -738
rect -1941 -772 -1925 -738
rect -1867 -772 -1851 -738
rect -1783 -772 -1767 -738
rect -1709 -772 -1693 -738
rect -1625 -772 -1609 -738
rect -1551 -772 -1535 -738
rect -1467 -772 -1451 -738
rect -1393 -772 -1377 -738
rect -1309 -772 -1293 -738
rect -1235 -772 -1219 -738
rect -1151 -772 -1135 -738
rect -1077 -772 -1061 -738
rect -993 -772 -977 -738
rect -919 -772 -903 -738
rect -835 -772 -819 -738
rect -761 -772 -745 -738
rect -677 -772 -661 -738
rect -603 -772 -587 -738
rect -519 -772 -503 -738
rect -445 -772 -429 -738
rect -361 -772 -345 -738
rect -287 -772 -271 -738
rect -203 -772 -187 -738
rect -129 -772 -113 -738
rect -45 -772 -29 -738
rect 29 -772 45 -738
rect 113 -772 129 -738
rect 187 -772 203 -738
rect 271 -772 287 -738
rect 345 -772 361 -738
rect 429 -772 445 -738
rect 503 -772 519 -738
rect 587 -772 603 -738
rect 661 -772 677 -738
rect 745 -772 761 -738
rect 819 -772 835 -738
rect 903 -772 919 -738
rect 977 -772 993 -738
rect 1061 -772 1077 -738
rect 1135 -772 1151 -738
rect 1219 -772 1235 -738
rect 1293 -772 1309 -738
rect 1377 -772 1393 -738
rect 1451 -772 1467 -738
rect 1535 -772 1551 -738
rect 1609 -772 1625 -738
rect 1693 -772 1709 -738
rect 1767 -772 1783 -738
rect 1851 -772 1867 -738
rect 1925 -772 1941 -738
rect 2009 -772 2025 -738
rect 2083 -772 2099 -738
rect 2167 -772 2183 -738
rect 2241 -772 2257 -738
rect 2325 -772 2341 -738
rect 2399 -772 2415 -738
rect 2483 -772 2499 -738
rect 2557 -772 2573 -738
rect 2641 -772 2657 -738
rect 2715 -772 2731 -738
rect 2799 -772 2815 -738
rect 2873 -772 2889 -738
rect 2957 -772 2973 -738
rect 3031 -772 3047 -738
rect 3115 -772 3131 -738
rect 3189 -772 3205 -738
rect 3273 -772 3289 -738
rect 3347 -772 3363 -738
rect 3431 -772 3447 -738
rect 3505 -772 3521 -738
rect 3589 -772 3605 -738
rect 3663 -772 3679 -738
rect 3747 -772 3763 -738
rect 3821 -772 3837 -738
rect 3905 -772 3921 -738
rect 3979 -772 3995 -738
rect 4063 -772 4079 -738
rect 4137 -772 4153 -738
rect 4221 -772 4237 -738
rect 4295 -772 4311 -738
rect 4379 -772 4395 -738
rect 4453 -772 4469 -738
rect 4537 -772 4553 -738
rect 4611 -772 4627 -738
rect 4695 -772 4711 -738
rect 4769 -772 4785 -738
rect 4853 -772 4869 -738
rect 4927 -772 4943 -738
rect 5011 -772 5027 -738
rect 5085 -772 5101 -738
rect 5169 -772 5185 -738
rect 5243 -772 5259 -738
rect 5327 -772 5343 -738
rect 5401 -772 5417 -738
rect 5485 -772 5501 -738
rect 5559 -772 5575 -738
rect 5643 -772 5659 -738
rect 5717 -772 5733 -738
rect 5801 -772 5817 -738
rect 5875 -772 5891 -738
rect 5959 -772 5975 -738
rect 6033 -772 6049 -738
rect 6117 -772 6133 -738
rect 6191 -772 6207 -738
rect 6275 -772 6291 -738
rect 6349 -772 6365 -738
rect 6433 -772 6449 -738
rect 6507 -772 6523 -738
rect 6591 -772 6607 -738
rect 6665 -772 6681 -738
rect 6749 -772 6765 -738
rect 6823 -772 6839 -738
rect 6907 -772 6923 -738
<< viali >>
rect -6969 -688 -6935 688
rect -6811 -688 -6777 688
rect -6653 -688 -6619 688
rect -6495 -688 -6461 688
rect -6337 -688 -6303 688
rect -6179 -688 -6145 688
rect -6021 -688 -5987 688
rect -5863 -688 -5829 688
rect -5705 -688 -5671 688
rect -5547 -688 -5513 688
rect -5389 -688 -5355 688
rect -5231 -688 -5197 688
rect -5073 -688 -5039 688
rect -4915 -688 -4881 688
rect -4757 -688 -4723 688
rect -4599 -688 -4565 688
rect -4441 -688 -4407 688
rect -4283 -688 -4249 688
rect -4125 -688 -4091 688
rect -3967 -688 -3933 688
rect -3809 -688 -3775 688
rect -3651 -688 -3617 688
rect -3493 -688 -3459 688
rect -3335 -688 -3301 688
rect -3177 -688 -3143 688
rect -3019 -688 -2985 688
rect -2861 -688 -2827 688
rect -2703 -688 -2669 688
rect -2545 -688 -2511 688
rect -2387 -688 -2353 688
rect -2229 -688 -2195 688
rect -2071 -688 -2037 688
rect -1913 -688 -1879 688
rect -1755 -688 -1721 688
rect -1597 -688 -1563 688
rect -1439 -688 -1405 688
rect -1281 -688 -1247 688
rect -1123 -688 -1089 688
rect -965 -688 -931 688
rect -807 -688 -773 688
rect -649 -688 -615 688
rect -491 -688 -457 688
rect -333 -688 -299 688
rect -175 -688 -141 688
rect -17 -688 17 688
rect 141 -688 175 688
rect 299 -688 333 688
rect 457 -688 491 688
rect 615 -688 649 688
rect 773 -688 807 688
rect 931 -688 965 688
rect 1089 -688 1123 688
rect 1247 -688 1281 688
rect 1405 -688 1439 688
rect 1563 -688 1597 688
rect 1721 -688 1755 688
rect 1879 -688 1913 688
rect 2037 -688 2071 688
rect 2195 -688 2229 688
rect 2353 -688 2387 688
rect 2511 -688 2545 688
rect 2669 -688 2703 688
rect 2827 -688 2861 688
rect 2985 -688 3019 688
rect 3143 -688 3177 688
rect 3301 -688 3335 688
rect 3459 -688 3493 688
rect 3617 -688 3651 688
rect 3775 -688 3809 688
rect 3933 -688 3967 688
rect 4091 -688 4125 688
rect 4249 -688 4283 688
rect 4407 -688 4441 688
rect 4565 -688 4599 688
rect 4723 -688 4757 688
rect 4881 -688 4915 688
rect 5039 -688 5073 688
rect 5197 -688 5231 688
rect 5355 -688 5389 688
rect 5513 -688 5547 688
rect 5671 -688 5705 688
rect 5829 -688 5863 688
rect 5987 -688 6021 688
rect 6145 -688 6179 688
rect 6303 -688 6337 688
rect 6461 -688 6495 688
rect 6619 -688 6653 688
rect 6777 -688 6811 688
rect 6935 -688 6969 688
<< metal1 >>
rect -6975 688 -6929 700
rect -6975 -688 -6969 688
rect -6935 -688 -6929 688
rect -6975 -700 -6929 -688
rect -6817 688 -6771 700
rect -6817 -688 -6811 688
rect -6777 -688 -6771 688
rect -6817 -700 -6771 -688
rect -6659 688 -6613 700
rect -6659 -688 -6653 688
rect -6619 -688 -6613 688
rect -6659 -700 -6613 -688
rect -6501 688 -6455 700
rect -6501 -688 -6495 688
rect -6461 -688 -6455 688
rect -6501 -700 -6455 -688
rect -6343 688 -6297 700
rect -6343 -688 -6337 688
rect -6303 -688 -6297 688
rect -6343 -700 -6297 -688
rect -6185 688 -6139 700
rect -6185 -688 -6179 688
rect -6145 -688 -6139 688
rect -6185 -700 -6139 -688
rect -6027 688 -5981 700
rect -6027 -688 -6021 688
rect -5987 -688 -5981 688
rect -6027 -700 -5981 -688
rect -5869 688 -5823 700
rect -5869 -688 -5863 688
rect -5829 -688 -5823 688
rect -5869 -700 -5823 -688
rect -5711 688 -5665 700
rect -5711 -688 -5705 688
rect -5671 -688 -5665 688
rect -5711 -700 -5665 -688
rect -5553 688 -5507 700
rect -5553 -688 -5547 688
rect -5513 -688 -5507 688
rect -5553 -700 -5507 -688
rect -5395 688 -5349 700
rect -5395 -688 -5389 688
rect -5355 -688 -5349 688
rect -5395 -700 -5349 -688
rect -5237 688 -5191 700
rect -5237 -688 -5231 688
rect -5197 -688 -5191 688
rect -5237 -700 -5191 -688
rect -5079 688 -5033 700
rect -5079 -688 -5073 688
rect -5039 -688 -5033 688
rect -5079 -700 -5033 -688
rect -4921 688 -4875 700
rect -4921 -688 -4915 688
rect -4881 -688 -4875 688
rect -4921 -700 -4875 -688
rect -4763 688 -4717 700
rect -4763 -688 -4757 688
rect -4723 -688 -4717 688
rect -4763 -700 -4717 -688
rect -4605 688 -4559 700
rect -4605 -688 -4599 688
rect -4565 -688 -4559 688
rect -4605 -700 -4559 -688
rect -4447 688 -4401 700
rect -4447 -688 -4441 688
rect -4407 -688 -4401 688
rect -4447 -700 -4401 -688
rect -4289 688 -4243 700
rect -4289 -688 -4283 688
rect -4249 -688 -4243 688
rect -4289 -700 -4243 -688
rect -4131 688 -4085 700
rect -4131 -688 -4125 688
rect -4091 -688 -4085 688
rect -4131 -700 -4085 -688
rect -3973 688 -3927 700
rect -3973 -688 -3967 688
rect -3933 -688 -3927 688
rect -3973 -700 -3927 -688
rect -3815 688 -3769 700
rect -3815 -688 -3809 688
rect -3775 -688 -3769 688
rect -3815 -700 -3769 -688
rect -3657 688 -3611 700
rect -3657 -688 -3651 688
rect -3617 -688 -3611 688
rect -3657 -700 -3611 -688
rect -3499 688 -3453 700
rect -3499 -688 -3493 688
rect -3459 -688 -3453 688
rect -3499 -700 -3453 -688
rect -3341 688 -3295 700
rect -3341 -688 -3335 688
rect -3301 -688 -3295 688
rect -3341 -700 -3295 -688
rect -3183 688 -3137 700
rect -3183 -688 -3177 688
rect -3143 -688 -3137 688
rect -3183 -700 -3137 -688
rect -3025 688 -2979 700
rect -3025 -688 -3019 688
rect -2985 -688 -2979 688
rect -3025 -700 -2979 -688
rect -2867 688 -2821 700
rect -2867 -688 -2861 688
rect -2827 -688 -2821 688
rect -2867 -700 -2821 -688
rect -2709 688 -2663 700
rect -2709 -688 -2703 688
rect -2669 -688 -2663 688
rect -2709 -700 -2663 -688
rect -2551 688 -2505 700
rect -2551 -688 -2545 688
rect -2511 -688 -2505 688
rect -2551 -700 -2505 -688
rect -2393 688 -2347 700
rect -2393 -688 -2387 688
rect -2353 -688 -2347 688
rect -2393 -700 -2347 -688
rect -2235 688 -2189 700
rect -2235 -688 -2229 688
rect -2195 -688 -2189 688
rect -2235 -700 -2189 -688
rect -2077 688 -2031 700
rect -2077 -688 -2071 688
rect -2037 -688 -2031 688
rect -2077 -700 -2031 -688
rect -1919 688 -1873 700
rect -1919 -688 -1913 688
rect -1879 -688 -1873 688
rect -1919 -700 -1873 -688
rect -1761 688 -1715 700
rect -1761 -688 -1755 688
rect -1721 -688 -1715 688
rect -1761 -700 -1715 -688
rect -1603 688 -1557 700
rect -1603 -688 -1597 688
rect -1563 -688 -1557 688
rect -1603 -700 -1557 -688
rect -1445 688 -1399 700
rect -1445 -688 -1439 688
rect -1405 -688 -1399 688
rect -1445 -700 -1399 -688
rect -1287 688 -1241 700
rect -1287 -688 -1281 688
rect -1247 -688 -1241 688
rect -1287 -700 -1241 -688
rect -1129 688 -1083 700
rect -1129 -688 -1123 688
rect -1089 -688 -1083 688
rect -1129 -700 -1083 -688
rect -971 688 -925 700
rect -971 -688 -965 688
rect -931 -688 -925 688
rect -971 -700 -925 -688
rect -813 688 -767 700
rect -813 -688 -807 688
rect -773 -688 -767 688
rect -813 -700 -767 -688
rect -655 688 -609 700
rect -655 -688 -649 688
rect -615 -688 -609 688
rect -655 -700 -609 -688
rect -497 688 -451 700
rect -497 -688 -491 688
rect -457 -688 -451 688
rect -497 -700 -451 -688
rect -339 688 -293 700
rect -339 -688 -333 688
rect -299 -688 -293 688
rect -339 -700 -293 -688
rect -181 688 -135 700
rect -181 -688 -175 688
rect -141 -688 -135 688
rect -181 -700 -135 -688
rect -23 688 23 700
rect -23 -688 -17 688
rect 17 -688 23 688
rect -23 -700 23 -688
rect 135 688 181 700
rect 135 -688 141 688
rect 175 -688 181 688
rect 135 -700 181 -688
rect 293 688 339 700
rect 293 -688 299 688
rect 333 -688 339 688
rect 293 -700 339 -688
rect 451 688 497 700
rect 451 -688 457 688
rect 491 -688 497 688
rect 451 -700 497 -688
rect 609 688 655 700
rect 609 -688 615 688
rect 649 -688 655 688
rect 609 -700 655 -688
rect 767 688 813 700
rect 767 -688 773 688
rect 807 -688 813 688
rect 767 -700 813 -688
rect 925 688 971 700
rect 925 -688 931 688
rect 965 -688 971 688
rect 925 -700 971 -688
rect 1083 688 1129 700
rect 1083 -688 1089 688
rect 1123 -688 1129 688
rect 1083 -700 1129 -688
rect 1241 688 1287 700
rect 1241 -688 1247 688
rect 1281 -688 1287 688
rect 1241 -700 1287 -688
rect 1399 688 1445 700
rect 1399 -688 1405 688
rect 1439 -688 1445 688
rect 1399 -700 1445 -688
rect 1557 688 1603 700
rect 1557 -688 1563 688
rect 1597 -688 1603 688
rect 1557 -700 1603 -688
rect 1715 688 1761 700
rect 1715 -688 1721 688
rect 1755 -688 1761 688
rect 1715 -700 1761 -688
rect 1873 688 1919 700
rect 1873 -688 1879 688
rect 1913 -688 1919 688
rect 1873 -700 1919 -688
rect 2031 688 2077 700
rect 2031 -688 2037 688
rect 2071 -688 2077 688
rect 2031 -700 2077 -688
rect 2189 688 2235 700
rect 2189 -688 2195 688
rect 2229 -688 2235 688
rect 2189 -700 2235 -688
rect 2347 688 2393 700
rect 2347 -688 2353 688
rect 2387 -688 2393 688
rect 2347 -700 2393 -688
rect 2505 688 2551 700
rect 2505 -688 2511 688
rect 2545 -688 2551 688
rect 2505 -700 2551 -688
rect 2663 688 2709 700
rect 2663 -688 2669 688
rect 2703 -688 2709 688
rect 2663 -700 2709 -688
rect 2821 688 2867 700
rect 2821 -688 2827 688
rect 2861 -688 2867 688
rect 2821 -700 2867 -688
rect 2979 688 3025 700
rect 2979 -688 2985 688
rect 3019 -688 3025 688
rect 2979 -700 3025 -688
rect 3137 688 3183 700
rect 3137 -688 3143 688
rect 3177 -688 3183 688
rect 3137 -700 3183 -688
rect 3295 688 3341 700
rect 3295 -688 3301 688
rect 3335 -688 3341 688
rect 3295 -700 3341 -688
rect 3453 688 3499 700
rect 3453 -688 3459 688
rect 3493 -688 3499 688
rect 3453 -700 3499 -688
rect 3611 688 3657 700
rect 3611 -688 3617 688
rect 3651 -688 3657 688
rect 3611 -700 3657 -688
rect 3769 688 3815 700
rect 3769 -688 3775 688
rect 3809 -688 3815 688
rect 3769 -700 3815 -688
rect 3927 688 3973 700
rect 3927 -688 3933 688
rect 3967 -688 3973 688
rect 3927 -700 3973 -688
rect 4085 688 4131 700
rect 4085 -688 4091 688
rect 4125 -688 4131 688
rect 4085 -700 4131 -688
rect 4243 688 4289 700
rect 4243 -688 4249 688
rect 4283 -688 4289 688
rect 4243 -700 4289 -688
rect 4401 688 4447 700
rect 4401 -688 4407 688
rect 4441 -688 4447 688
rect 4401 -700 4447 -688
rect 4559 688 4605 700
rect 4559 -688 4565 688
rect 4599 -688 4605 688
rect 4559 -700 4605 -688
rect 4717 688 4763 700
rect 4717 -688 4723 688
rect 4757 -688 4763 688
rect 4717 -700 4763 -688
rect 4875 688 4921 700
rect 4875 -688 4881 688
rect 4915 -688 4921 688
rect 4875 -700 4921 -688
rect 5033 688 5079 700
rect 5033 -688 5039 688
rect 5073 -688 5079 688
rect 5033 -700 5079 -688
rect 5191 688 5237 700
rect 5191 -688 5197 688
rect 5231 -688 5237 688
rect 5191 -700 5237 -688
rect 5349 688 5395 700
rect 5349 -688 5355 688
rect 5389 -688 5395 688
rect 5349 -700 5395 -688
rect 5507 688 5553 700
rect 5507 -688 5513 688
rect 5547 -688 5553 688
rect 5507 -700 5553 -688
rect 5665 688 5711 700
rect 5665 -688 5671 688
rect 5705 -688 5711 688
rect 5665 -700 5711 -688
rect 5823 688 5869 700
rect 5823 -688 5829 688
rect 5863 -688 5869 688
rect 5823 -700 5869 -688
rect 5981 688 6027 700
rect 5981 -688 5987 688
rect 6021 -688 6027 688
rect 5981 -700 6027 -688
rect 6139 688 6185 700
rect 6139 -688 6145 688
rect 6179 -688 6185 688
rect 6139 -700 6185 -688
rect 6297 688 6343 700
rect 6297 -688 6303 688
rect 6337 -688 6343 688
rect 6297 -700 6343 -688
rect 6455 688 6501 700
rect 6455 -688 6461 688
rect 6495 -688 6501 688
rect 6455 -700 6501 -688
rect 6613 688 6659 700
rect 6613 -688 6619 688
rect 6653 -688 6659 688
rect 6613 -700 6659 -688
rect 6771 688 6817 700
rect 6771 -688 6777 688
rect 6811 -688 6817 688
rect 6771 -700 6817 -688
rect 6929 688 6975 700
rect 6929 -688 6935 688
rect 6969 -688 6975 688
rect 6929 -700 6975 -688
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 7 l 0.5 m 1 nf 88 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
