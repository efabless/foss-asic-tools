magic
tech sky130A
magscale 1 2
timestamp 1621030523
<< mvnmos >>
rect -100 -500 100 500
<< mvndiff >>
rect -158 488 -100 500
rect -158 -488 -146 488
rect -112 -488 -100 488
rect -158 -500 -100 -488
rect 100 488 158 500
rect 100 -488 112 488
rect 146 -488 158 488
rect 100 -500 158 -488
<< mvndiffc >>
rect -146 -488 -112 488
rect 112 -488 146 488
<< poly >>
rect -66 572 66 588
rect -66 555 -50 572
rect -100 538 -50 555
rect 50 555 66 572
rect 50 538 100 555
rect -100 500 100 538
rect -100 -538 100 -500
rect -100 -555 -50 -538
rect -66 -572 -50 -555
rect 50 -555 100 -538
rect 50 -572 66 -555
rect -66 -588 66 -572
<< polycont >>
rect -50 538 50 572
rect -50 -572 50 -538
<< locali >>
rect -66 538 -50 572
rect 50 538 66 572
rect -146 488 -112 504
rect -146 -504 -112 -488
rect 112 488 146 504
rect 112 -504 146 -488
rect -66 -572 -50 -538
rect 50 -572 66 -538
<< viali >>
rect -34 538 34 572
rect -146 -488 -112 488
rect 112 -488 146 488
rect -34 -572 34 -538
<< metal1 >>
rect -46 572 46 578
rect -46 538 -34 572
rect 34 538 46 572
rect -46 532 46 538
rect -152 488 -106 500
rect -152 -488 -146 488
rect -112 -488 -106 488
rect -152 -500 -106 -488
rect 106 488 152 500
rect 106 -488 112 488
rect 146 -488 152 488
rect 106 -500 152 -488
rect -46 -538 46 -532
rect -46 -572 -34 -538
rect 34 -572 46 -538
rect -46 -578 46 -572
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 5 l 1 m 1 nf 1 diffcov 100 polycov 60 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
