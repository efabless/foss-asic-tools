magic
tech sky130A
timestamp 1384693831
<< checkpaint >>
rect -630 -615 888 2142
use INV_28319830_0_0_1678192857  INV_28319830_0_0_1678192857_0
timestamp 1384693831
transform 1 0 0 0 1 0
box 0 15 258 1512
<< labels >>
flabel metal1 s 172 294 172 294 0 FreeSerif 0 0 0 0 A
flabel metal2 s 86 378 86 378 0 FreeSerif 0 0 0 0 VSS
flabel metal2 s 86 1134 86 1134 0 FreeSerif 0 0 0 0 VDD
flabel metal1 s 172 714 172 714 0 FreeSerif 0 0 0 0 Y
<< end >>
