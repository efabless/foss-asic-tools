magic
tech sky130A
magscale 1 2
timestamp 1620937039
<< error_p >>
rect -224 -566 -194 566
rect -158 -500 -128 500
rect 128 -500 158 500
rect 194 -566 224 566
<< nwell >>
rect -194 -600 194 600
<< mvpmos >>
rect -100 -500 100 500
<< mvpdiff >>
rect -158 488 -100 500
rect -158 -488 -146 488
rect -112 -488 -100 488
rect -158 -500 -100 -488
rect 100 488 158 500
rect 100 -488 112 488
rect 146 -488 158 488
rect 100 -500 158 -488
<< mvpdiffc >>
rect -146 -488 -112 488
rect 112 -488 146 488
<< poly >>
rect -66 581 66 597
rect -66 564 -50 581
rect -100 547 -50 564
rect 50 564 66 581
rect 50 547 100 564
rect -100 500 100 547
rect -100 -547 100 -500
rect -100 -564 -50 -547
rect -66 -581 -50 -564
rect 50 -564 100 -547
rect 50 -581 66 -564
rect -66 -597 66 -581
<< polycont >>
rect -50 547 50 581
rect -50 -581 50 -547
<< locali >>
rect -66 547 -50 581
rect 50 547 66 581
rect -146 488 -112 504
rect -146 -504 -112 -488
rect 112 488 146 504
rect 112 -504 146 -488
rect -66 -581 -50 -547
rect 50 -581 66 -547
<< viali >>
rect -34 547 34 581
rect -146 -488 -112 488
rect 112 -488 146 488
rect -34 -581 34 -547
<< metal1 >>
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect -152 488 -106 500
rect -152 -488 -146 488
rect -112 -488 -106 488
rect -152 -500 -106 -488
rect 106 488 152 500
rect 106 -488 112 488
rect 146 -488 152 488
rect 106 -500 152 -488
rect -46 -547 46 -541
rect -46 -581 -34 -547
rect 34 -581 46 -547
rect -46 -587 46 -581
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 5 l 1 m 1 nf 1 diffcov 100 polycov 60 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
