magic
tech sky130A
magscale 1 2
timestamp 1624430562
<< error_p >>
rect -2129 566 2129 600
rect -2159 -566 2159 566
rect -2129 -600 2129 -566
<< nwell >>
rect -2129 -600 2129 600
<< mvpmos >>
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
<< mvpdiff >>
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
<< mvpdiffc >>
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
<< poly >>
rect -2001 581 -1869 597
rect -2001 564 -1985 581
rect -2035 547 -1985 564
rect -1885 564 -1869 581
rect -1743 581 -1611 597
rect -1743 564 -1727 581
rect -1885 547 -1835 564
rect -2035 500 -1835 547
rect -1777 547 -1727 564
rect -1627 564 -1611 581
rect -1485 581 -1353 597
rect -1485 564 -1469 581
rect -1627 547 -1577 564
rect -1777 500 -1577 547
rect -1519 547 -1469 564
rect -1369 564 -1353 581
rect -1227 581 -1095 597
rect -1227 564 -1211 581
rect -1369 547 -1319 564
rect -1519 500 -1319 547
rect -1261 547 -1211 564
rect -1111 564 -1095 581
rect -969 581 -837 597
rect -969 564 -953 581
rect -1111 547 -1061 564
rect -1261 500 -1061 547
rect -1003 547 -953 564
rect -853 564 -837 581
rect -711 581 -579 597
rect -711 564 -695 581
rect -853 547 -803 564
rect -1003 500 -803 547
rect -745 547 -695 564
rect -595 564 -579 581
rect -453 581 -321 597
rect -453 564 -437 581
rect -595 547 -545 564
rect -745 500 -545 547
rect -487 547 -437 564
rect -337 564 -321 581
rect -195 581 -63 597
rect -195 564 -179 581
rect -337 547 -287 564
rect -487 500 -287 547
rect -229 547 -179 564
rect -79 564 -63 581
rect 63 581 195 597
rect 63 564 79 581
rect -79 547 -29 564
rect -229 500 -29 547
rect 29 547 79 564
rect 179 564 195 581
rect 321 581 453 597
rect 321 564 337 581
rect 179 547 229 564
rect 29 500 229 547
rect 287 547 337 564
rect 437 564 453 581
rect 579 581 711 597
rect 579 564 595 581
rect 437 547 487 564
rect 287 500 487 547
rect 545 547 595 564
rect 695 564 711 581
rect 837 581 969 597
rect 837 564 853 581
rect 695 547 745 564
rect 545 500 745 547
rect 803 547 853 564
rect 953 564 969 581
rect 1095 581 1227 597
rect 1095 564 1111 581
rect 953 547 1003 564
rect 803 500 1003 547
rect 1061 547 1111 564
rect 1211 564 1227 581
rect 1353 581 1485 597
rect 1353 564 1369 581
rect 1211 547 1261 564
rect 1061 500 1261 547
rect 1319 547 1369 564
rect 1469 564 1485 581
rect 1611 581 1743 597
rect 1611 564 1627 581
rect 1469 547 1519 564
rect 1319 500 1519 547
rect 1577 547 1627 564
rect 1727 564 1743 581
rect 1869 581 2001 597
rect 1869 564 1885 581
rect 1727 547 1777 564
rect 1577 500 1777 547
rect 1835 547 1885 564
rect 1985 564 2001 581
rect 1985 547 2035 564
rect 1835 500 2035 547
rect -2035 -547 -1835 -500
rect -2035 -564 -1985 -547
rect -2001 -581 -1985 -564
rect -1885 -564 -1835 -547
rect -1777 -547 -1577 -500
rect -1777 -564 -1727 -547
rect -1885 -581 -1869 -564
rect -2001 -597 -1869 -581
rect -1743 -581 -1727 -564
rect -1627 -564 -1577 -547
rect -1519 -547 -1319 -500
rect -1519 -564 -1469 -547
rect -1627 -581 -1611 -564
rect -1743 -597 -1611 -581
rect -1485 -581 -1469 -564
rect -1369 -564 -1319 -547
rect -1261 -547 -1061 -500
rect -1261 -564 -1211 -547
rect -1369 -581 -1353 -564
rect -1485 -597 -1353 -581
rect -1227 -581 -1211 -564
rect -1111 -564 -1061 -547
rect -1003 -547 -803 -500
rect -1003 -564 -953 -547
rect -1111 -581 -1095 -564
rect -1227 -597 -1095 -581
rect -969 -581 -953 -564
rect -853 -564 -803 -547
rect -745 -547 -545 -500
rect -745 -564 -695 -547
rect -853 -581 -837 -564
rect -969 -597 -837 -581
rect -711 -581 -695 -564
rect -595 -564 -545 -547
rect -487 -547 -287 -500
rect -487 -564 -437 -547
rect -595 -581 -579 -564
rect -711 -597 -579 -581
rect -453 -581 -437 -564
rect -337 -564 -287 -547
rect -229 -547 -29 -500
rect -229 -564 -179 -547
rect -337 -581 -321 -564
rect -453 -597 -321 -581
rect -195 -581 -179 -564
rect -79 -564 -29 -547
rect 29 -547 229 -500
rect 29 -564 79 -547
rect -79 -581 -63 -564
rect -195 -597 -63 -581
rect 63 -581 79 -564
rect 179 -564 229 -547
rect 287 -547 487 -500
rect 287 -564 337 -547
rect 179 -581 195 -564
rect 63 -597 195 -581
rect 321 -581 337 -564
rect 437 -564 487 -547
rect 545 -547 745 -500
rect 545 -564 595 -547
rect 437 -581 453 -564
rect 321 -597 453 -581
rect 579 -581 595 -564
rect 695 -564 745 -547
rect 803 -547 1003 -500
rect 803 -564 853 -547
rect 695 -581 711 -564
rect 579 -597 711 -581
rect 837 -581 853 -564
rect 953 -564 1003 -547
rect 1061 -547 1261 -500
rect 1061 -564 1111 -547
rect 953 -581 969 -564
rect 837 -597 969 -581
rect 1095 -581 1111 -564
rect 1211 -564 1261 -547
rect 1319 -547 1519 -500
rect 1319 -564 1369 -547
rect 1211 -581 1227 -564
rect 1095 -597 1227 -581
rect 1353 -581 1369 -564
rect 1469 -564 1519 -547
rect 1577 -547 1777 -500
rect 1577 -564 1627 -547
rect 1469 -581 1485 -564
rect 1353 -597 1485 -581
rect 1611 -581 1627 -564
rect 1727 -564 1777 -547
rect 1835 -547 2035 -500
rect 1835 -564 1885 -547
rect 1727 -581 1743 -564
rect 1611 -597 1743 -581
rect 1869 -581 1885 -564
rect 1985 -564 2035 -547
rect 1985 -581 2001 -564
rect 1869 -597 2001 -581
<< polycont >>
rect -1985 547 -1885 581
rect -1727 547 -1627 581
rect -1469 547 -1369 581
rect -1211 547 -1111 581
rect -953 547 -853 581
rect -695 547 -595 581
rect -437 547 -337 581
rect -179 547 -79 581
rect 79 547 179 581
rect 337 547 437 581
rect 595 547 695 581
rect 853 547 953 581
rect 1111 547 1211 581
rect 1369 547 1469 581
rect 1627 547 1727 581
rect 1885 547 1985 581
rect -1985 -581 -1885 -547
rect -1727 -581 -1627 -547
rect -1469 -581 -1369 -547
rect -1211 -581 -1111 -547
rect -953 -581 -853 -547
rect -695 -581 -595 -547
rect -437 -581 -337 -547
rect -179 -581 -79 -547
rect 79 -581 179 -547
rect 337 -581 437 -547
rect 595 -581 695 -547
rect 853 -581 953 -547
rect 1111 -581 1211 -547
rect 1369 -581 1469 -547
rect 1627 -581 1727 -547
rect 1885 -581 1985 -547
<< locali >>
rect -2001 547 -1985 581
rect -1885 547 -1869 581
rect -1743 547 -1727 581
rect -1627 547 -1611 581
rect -1485 547 -1469 581
rect -1369 547 -1353 581
rect -1227 547 -1211 581
rect -1111 547 -1095 581
rect -969 547 -953 581
rect -853 547 -837 581
rect -711 547 -695 581
rect -595 547 -579 581
rect -453 547 -437 581
rect -337 547 -321 581
rect -195 547 -179 581
rect -79 547 -63 581
rect 63 547 79 581
rect 179 547 195 581
rect 321 547 337 581
rect 437 547 453 581
rect 579 547 595 581
rect 695 547 711 581
rect 837 547 853 581
rect 953 547 969 581
rect 1095 547 1111 581
rect 1211 547 1227 581
rect 1353 547 1369 581
rect 1469 547 1485 581
rect 1611 547 1627 581
rect 1727 547 1743 581
rect 1869 547 1885 581
rect 1985 547 2001 581
rect -2081 488 -2047 504
rect -2081 -504 -2047 -488
rect -1823 488 -1789 504
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect 1789 488 1823 504
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -504 2081 -488
rect -2001 -581 -1985 -547
rect -1885 -581 -1869 -547
rect -1743 -581 -1727 -547
rect -1627 -581 -1611 -547
rect -1485 -581 -1469 -547
rect -1369 -581 -1353 -547
rect -1227 -581 -1211 -547
rect -1111 -581 -1095 -547
rect -969 -581 -953 -547
rect -853 -581 -837 -547
rect -711 -581 -695 -547
rect -595 -581 -579 -547
rect -453 -581 -437 -547
rect -337 -581 -321 -547
rect -195 -581 -179 -547
rect -79 -581 -63 -547
rect 63 -581 79 -547
rect 179 -581 195 -547
rect 321 -581 337 -547
rect 437 -581 453 -547
rect 579 -581 595 -547
rect 695 -581 711 -547
rect 837 -581 853 -547
rect 953 -581 969 -547
rect 1095 -581 1111 -547
rect 1211 -581 1227 -547
rect 1353 -581 1369 -547
rect 1469 -581 1485 -547
rect 1611 -581 1627 -547
rect 1727 -581 1743 -547
rect 1869 -581 1885 -547
rect 1985 -581 2001 -547
<< viali >>
rect -1969 547 -1901 581
rect -1711 547 -1643 581
rect -1453 547 -1385 581
rect -1195 547 -1127 581
rect -937 547 -869 581
rect -679 547 -611 581
rect -421 547 -353 581
rect -163 547 -95 581
rect 95 547 163 581
rect 353 547 421 581
rect 611 547 679 581
rect 869 547 937 581
rect 1127 547 1195 581
rect 1385 547 1453 581
rect 1643 547 1711 581
rect 1901 547 1969 581
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect -1969 -581 -1901 -547
rect -1711 -581 -1643 -547
rect -1453 -581 -1385 -547
rect -1195 -581 -1127 -547
rect -937 -581 -869 -547
rect -679 -581 -611 -547
rect -421 -581 -353 -547
rect -163 -581 -95 -547
rect 95 -581 163 -547
rect 353 -581 421 -547
rect 611 -581 679 -547
rect 869 -581 937 -547
rect 1127 -581 1195 -547
rect 1385 -581 1453 -547
rect 1643 -581 1711 -547
rect 1901 -581 1969 -547
<< metal1 >>
rect -1981 581 -1889 587
rect -1981 547 -1969 581
rect -1901 547 -1889 581
rect -1981 541 -1889 547
rect -1723 581 -1631 587
rect -1723 547 -1711 581
rect -1643 547 -1631 581
rect -1723 541 -1631 547
rect -1465 581 -1373 587
rect -1465 547 -1453 581
rect -1385 547 -1373 581
rect -1465 541 -1373 547
rect -1207 581 -1115 587
rect -1207 547 -1195 581
rect -1127 547 -1115 581
rect -1207 541 -1115 547
rect -949 581 -857 587
rect -949 547 -937 581
rect -869 547 -857 581
rect -949 541 -857 547
rect -691 581 -599 587
rect -691 547 -679 581
rect -611 547 -599 581
rect -691 541 -599 547
rect -433 581 -341 587
rect -433 547 -421 581
rect -353 547 -341 581
rect -433 541 -341 547
rect -175 581 -83 587
rect -175 547 -163 581
rect -95 547 -83 581
rect -175 541 -83 547
rect 83 581 175 587
rect 83 547 95 581
rect 163 547 175 581
rect 83 541 175 547
rect 341 581 433 587
rect 341 547 353 581
rect 421 547 433 581
rect 341 541 433 547
rect 599 581 691 587
rect 599 547 611 581
rect 679 547 691 581
rect 599 541 691 547
rect 857 581 949 587
rect 857 547 869 581
rect 937 547 949 581
rect 857 541 949 547
rect 1115 581 1207 587
rect 1115 547 1127 581
rect 1195 547 1207 581
rect 1115 541 1207 547
rect 1373 581 1465 587
rect 1373 547 1385 581
rect 1453 547 1465 581
rect 1373 541 1465 547
rect 1631 581 1723 587
rect 1631 547 1643 581
rect 1711 547 1723 581
rect 1631 541 1723 547
rect 1889 581 1981 587
rect 1889 547 1901 581
rect 1969 547 1981 581
rect 1889 541 1981 547
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
rect -1981 -547 -1889 -541
rect -1981 -581 -1969 -547
rect -1901 -581 -1889 -547
rect -1981 -587 -1889 -581
rect -1723 -547 -1631 -541
rect -1723 -581 -1711 -547
rect -1643 -581 -1631 -547
rect -1723 -587 -1631 -581
rect -1465 -547 -1373 -541
rect -1465 -581 -1453 -547
rect -1385 -581 -1373 -547
rect -1465 -587 -1373 -581
rect -1207 -547 -1115 -541
rect -1207 -581 -1195 -547
rect -1127 -581 -1115 -547
rect -1207 -587 -1115 -581
rect -949 -547 -857 -541
rect -949 -581 -937 -547
rect -869 -581 -857 -547
rect -949 -587 -857 -581
rect -691 -547 -599 -541
rect -691 -581 -679 -547
rect -611 -581 -599 -547
rect -691 -587 -599 -581
rect -433 -547 -341 -541
rect -433 -581 -421 -547
rect -353 -581 -341 -547
rect -433 -587 -341 -581
rect -175 -547 -83 -541
rect -175 -581 -163 -547
rect -95 -581 -83 -547
rect -175 -587 -83 -581
rect 83 -547 175 -541
rect 83 -581 95 -547
rect 163 -581 175 -547
rect 83 -587 175 -581
rect 341 -547 433 -541
rect 341 -581 353 -547
rect 421 -581 433 -547
rect 341 -587 433 -581
rect 599 -547 691 -541
rect 599 -581 611 -547
rect 679 -581 691 -547
rect 599 -587 691 -581
rect 857 -547 949 -541
rect 857 -581 869 -547
rect 937 -581 949 -547
rect 857 -587 949 -581
rect 1115 -547 1207 -541
rect 1115 -581 1127 -547
rect 1195 -581 1207 -547
rect 1115 -587 1207 -581
rect 1373 -547 1465 -541
rect 1373 -581 1385 -547
rect 1453 -581 1465 -547
rect 1373 -587 1465 -581
rect 1631 -547 1723 -541
rect 1631 -581 1643 -547
rect 1711 -581 1723 -547
rect 1631 -587 1723 -581
rect 1889 -547 1981 -541
rect 1889 -581 1901 -547
rect 1969 -581 1981 -547
rect 1889 -587 1981 -581
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 5 l 1 m 1 nf 16 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
