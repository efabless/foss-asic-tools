magic
tech sky130A
magscale 1 2
timestamp 1621838304
<< nwell >>
rect -3000 40 3000 4500
<< pwell >>
rect -3000 -4500 3000 -40
<< mvnmos >>
rect -1677 -1700 -1477 -700
rect -1419 -1700 -1319 -700
rect 1319 -1700 1419 -700
rect 1477 -1700 1677 -700
<< mvpmos >>
rect -1677 700 -1477 1700
rect -1419 700 -1319 1700
rect 1319 700 1419 1700
rect 1477 700 1677 1700
<< mvndiff >>
rect -1735 -712 -1677 -700
rect -1735 -1688 -1723 -712
rect -1689 -1688 -1677 -712
rect -1735 -1700 -1677 -1688
rect -1477 -712 -1419 -700
rect -1477 -1688 -1465 -712
rect -1431 -1688 -1419 -712
rect -1477 -1700 -1419 -1688
rect 1419 -712 1477 -700
rect 1419 -1688 1431 -712
rect 1465 -1688 1477 -712
rect 1419 -1700 1477 -1688
rect 1677 -712 1735 -700
rect 1677 -1688 1689 -712
rect 1723 -1688 1735 -712
rect 1677 -1700 1735 -1688
<< mvpdiff >>
rect -1735 1688 -1677 1700
rect -1735 712 -1723 1688
rect -1689 712 -1677 1688
rect -1735 700 -1677 712
rect -1477 1688 -1419 1700
rect -1477 712 -1465 1688
rect -1431 712 -1419 1688
rect -1477 700 -1419 712
rect 1419 1688 1477 1700
rect 1419 712 1431 1688
rect 1465 712 1477 1688
rect 1419 700 1477 712
rect 1677 1688 1735 1700
rect 1677 712 1689 1688
rect 1723 712 1735 1688
rect 1677 700 1735 712
<< mvndiffc >>
rect -1723 -1688 -1689 -712
rect -1465 -1688 -1431 -712
rect 1431 -1688 1465 -712
rect 1689 -1688 1723 -712
<< mvpdiffc >>
rect -1723 712 -1689 1688
rect -1465 712 -1431 1688
rect 1431 712 1465 1688
rect 1689 712 1723 1688
<< mvpsubdiff >>
rect -2934 -118 2934 -106
rect -2934 -218 -2760 -118
rect 2760 -218 2934 -118
rect -2934 -230 2934 -218
rect -2934 -280 -2810 -230
rect -2934 -4260 -2922 -280
rect -2822 -4260 -2810 -280
rect 2810 -280 2934 -230
rect -2934 -4310 -2810 -4260
rect 2810 -4260 2822 -280
rect 2922 -4260 2934 -280
rect 2810 -4310 2934 -4260
rect -2934 -4322 2934 -4310
rect -2934 -4422 -2760 -4322
rect 2760 -4422 2934 -4322
rect -2934 -4434 2934 -4422
<< mvnsubdiff >>
rect -2934 4422 2934 4434
rect -2934 4322 -2760 4422
rect 2760 4322 2934 4422
rect -2934 4310 2934 4322
rect -2934 4260 -2810 4310
rect -2934 280 -2922 4260
rect -2822 280 -2810 4260
rect 2810 4260 2934 4310
rect -2934 230 -2810 280
rect 2810 280 2822 4260
rect 2922 280 2934 4260
rect 2810 230 2934 280
rect -2934 218 2934 230
rect -2934 118 -2760 218
rect 2760 118 2934 218
rect -2934 106 2934 118
<< mvpsubdiffcont >>
rect -2760 -218 2760 -118
rect -2922 -4260 -2822 -280
rect 2822 -4260 2922 -280
rect -2760 -4422 2760 -4322
<< mvnsubdiffcont >>
rect -2760 4322 2760 4422
rect -2922 280 -2822 4260
rect 2822 280 2922 4260
rect -2760 118 2760 218
<< poly >>
rect -1643 1781 -1511 1797
rect -1643 1764 -1627 1781
rect -1677 1747 -1627 1764
rect -1527 1764 -1511 1781
rect -1419 1781 -1319 1797
rect -1527 1747 -1477 1764
rect -1677 1700 -1477 1747
rect -1419 1747 -1403 1781
rect -1335 1747 -1319 1781
rect -1419 1700 -1319 1747
rect -1677 653 -1477 700
rect -1677 636 -1627 653
rect -1643 619 -1627 636
rect -1527 636 -1477 653
rect -1419 653 -1319 700
rect -1527 619 -1511 636
rect -1643 603 -1511 619
rect -1419 619 -1403 653
rect -1335 619 -1319 653
rect -1419 603 -1319 619
rect 1319 1781 1419 1797
rect 1319 1747 1335 1781
rect 1403 1747 1419 1781
rect 1511 1781 1643 1797
rect 1511 1764 1527 1781
rect 1319 1700 1419 1747
rect 1477 1747 1527 1764
rect 1627 1764 1643 1781
rect 1627 1747 1677 1764
rect 1477 1700 1677 1747
rect 1319 653 1419 700
rect 1319 619 1335 653
rect 1403 619 1419 653
rect 1477 653 1677 700
rect 1477 636 1527 653
rect 1319 603 1419 619
rect 1511 619 1527 636
rect 1627 636 1677 653
rect 1627 619 1643 636
rect 1511 603 1643 619
rect -1643 -628 -1511 -612
rect -1643 -645 -1627 -628
rect -1677 -662 -1627 -645
rect -1527 -645 -1511 -628
rect -1419 -628 -1319 -612
rect -1527 -662 -1477 -645
rect -1677 -700 -1477 -662
rect -1419 -662 -1403 -628
rect -1335 -662 -1319 -628
rect -1419 -700 -1319 -662
rect -1677 -1738 -1477 -1700
rect -1677 -1755 -1627 -1738
rect -1643 -1772 -1627 -1755
rect -1527 -1755 -1477 -1738
rect -1419 -1738 -1319 -1700
rect -1527 -1772 -1511 -1755
rect -1643 -1788 -1511 -1772
rect -1419 -1772 -1403 -1738
rect -1335 -1772 -1319 -1738
rect -1419 -1788 -1319 -1772
rect 1319 -628 1419 -612
rect 1319 -662 1335 -628
rect 1403 -662 1419 -628
rect 1511 -628 1643 -612
rect 1511 -645 1527 -628
rect 1319 -700 1419 -662
rect 1477 -662 1527 -645
rect 1627 -645 1643 -628
rect 1627 -662 1677 -645
rect 1477 -700 1677 -662
rect 1319 -1738 1419 -1700
rect 1319 -1772 1335 -1738
rect 1403 -1772 1419 -1738
rect 1477 -1738 1677 -1700
rect 1477 -1755 1527 -1738
rect 1319 -1788 1419 -1772
rect 1511 -1772 1527 -1755
rect 1627 -1755 1677 -1738
rect 1627 -1772 1643 -1755
rect 1511 -1788 1643 -1772
<< polycont >>
rect -1627 1747 -1527 1781
rect -1403 1747 -1335 1781
rect -1627 619 -1527 653
rect -1403 619 -1335 653
rect 1335 1747 1403 1781
rect 1527 1747 1627 1781
rect 1335 619 1403 653
rect 1527 619 1627 653
rect -1627 -662 -1527 -628
rect -1403 -662 -1335 -628
rect -1627 -1772 -1527 -1738
rect -1403 -1772 -1335 -1738
rect 1335 -662 1403 -628
rect 1527 -662 1627 -628
rect 1335 -1772 1403 -1738
rect 1527 -1772 1627 -1738
<< locali >>
rect -2922 4260 -2822 4422
rect 2822 4260 2922 4422
rect -2001 3797 2001 4197
rect -2001 3547 -1869 3797
rect -1743 3547 -1611 3797
rect -1485 3547 -1353 3797
rect -969 3547 -837 3797
rect -711 3621 711 3763
rect -711 3547 -579 3621
rect -453 3547 -321 3621
rect -195 3547 -63 3621
rect 62 3547 195 3621
rect 321 3547 453 3621
rect 579 3547 711 3621
rect 837 3547 969 3797
rect 1353 3547 1485 3797
rect 1611 3547 1743 3797
rect 1869 3547 2001 3797
rect -1419 2282 1419 2333
rect -1419 2202 -659 2282
rect -579 2202 579 2282
rect 659 2202 1419 2282
rect -1419 2049 1419 2202
rect -1419 1781 -1319 2049
rect -1643 1747 -1627 1781
rect -1527 1747 -1511 1781
rect -1419 1747 -1403 1781
rect -1335 1747 -1319 1781
rect -969 2008 969 2015
rect -969 1958 -963 2008
rect -913 1958 913 2008
rect 963 1958 969 2008
rect -969 1821 969 1958
rect -969 1747 -837 1821
rect -195 1747 -63 1821
rect 63 1747 195 1821
rect 837 1747 969 1821
rect 1319 1781 1419 2049
rect 1319 1747 1335 1781
rect 1403 1747 1419 1781
rect 1511 1747 1527 1781
rect 1627 1747 1643 1781
rect -1723 1688 -1689 1704
rect -1723 696 -1689 712
rect -1465 1688 -1431 1704
rect -1465 696 -1431 712
rect 1431 1688 1465 1704
rect 1431 696 1465 712
rect 1689 1688 1723 1704
rect 1689 696 1723 712
rect -1643 619 -1627 653
rect -1527 619 -1511 653
rect -1419 619 -1403 653
rect -1335 619 -1319 653
rect -711 579 -579 653
rect -453 579 -321 653
rect 321 579 453 653
rect 579 579 711 653
rect 1319 619 1335 653
rect 1403 619 1419 653
rect 1511 619 1527 653
rect 1627 619 1643 653
rect -1262 567 1264 579
rect -1212 517 1202 567
rect 1252 517 1264 567
rect -1262 437 1264 517
rect -447 436 -315 437
rect -2922 118 -2822 280
rect 2822 118 2922 280
rect -2922 -280 -2822 -118
rect 2822 -280 2922 -118
rect -969 -458 969 -394
rect -969 -538 -41 -458
rect 39 -538 969 -458
rect -969 -588 969 -538
rect -1643 -662 -1627 -628
rect -1527 -662 -1511 -628
rect -1419 -662 -1403 -628
rect -1335 -662 -1319 -628
rect -969 -662 -837 -588
rect -195 -662 -63 -588
rect 63 -662 195 -588
rect 837 -662 969 -588
rect 1319 -662 1335 -628
rect 1403 -662 1419 -628
rect 1511 -662 1527 -628
rect 1627 -662 1643 -628
rect -1723 -712 -1689 -696
rect -1723 -1704 -1689 -1688
rect -1465 -712 -1431 -696
rect -1465 -1704 -1431 -1688
rect 1431 -712 1465 -696
rect 1431 -1704 1465 -1688
rect 1689 -712 1723 -696
rect 1689 -1704 1723 -1688
rect -1643 -1772 -1627 -1738
rect -1527 -1772 -1511 -1738
rect -1419 -1772 -1403 -1738
rect -1335 -1772 -1319 -1738
rect -1419 -1988 -1319 -1772
rect -711 -1812 -579 -1738
rect -453 -1812 -321 -1738
rect 321 -1812 453 -1738
rect 579 -1812 711 -1738
rect -711 -1822 711 -1812
rect -711 -1902 -685 -1822
rect -605 -1902 -427 -1822
rect -347 -1902 347 -1822
rect 427 -1902 605 -1822
rect 685 -1902 711 -1822
rect -711 -1954 711 -1902
rect 1319 -1772 1335 -1738
rect 1403 -1772 1419 -1738
rect 1511 -1772 1527 -1738
rect 1627 -1772 1643 -1738
rect 1319 -1988 1419 -1772
rect -1419 -2046 1419 -1988
rect -1419 -2126 -556 -2046
rect -476 -2126 476 -2046
rect 556 -2126 1419 -2046
rect -1419 -2272 1419 -2126
rect -2922 -4422 -2822 -4260
rect 2822 -4422 2922 -4260
<< viali >>
rect -2822 4322 -2760 4422
rect -2760 4322 2760 4422
rect 2760 4322 2822 4422
rect -2922 423 -2822 4117
rect -659 2202 -579 2282
rect 579 2202 659 2282
rect -1611 1747 -1543 1781
rect -1396 1747 -1342 1781
rect -963 1958 -913 2008
rect 913 1958 963 2008
rect 1342 1747 1396 1781
rect 1543 1747 1611 1781
rect -1723 712 -1689 1688
rect -1465 712 -1431 1688
rect 1431 712 1465 1688
rect 1689 712 1723 1688
rect -1611 619 -1543 653
rect -1396 619 -1342 653
rect 1342 619 1396 653
rect 1543 619 1611 653
rect -1262 517 -1212 567
rect 1202 517 1252 567
rect 2822 423 2922 4117
rect -2822 118 -2760 218
rect -2760 118 2760 218
rect 2760 118 2822 218
rect -2822 -218 -2760 -118
rect -2760 -218 2760 -118
rect 2760 -218 2822 -118
rect -2922 -4117 -2822 -423
rect -41 -538 39 -458
rect -1611 -662 -1543 -628
rect -1396 -662 -1342 -628
rect 1342 -662 1396 -628
rect 1543 -662 1611 -628
rect -1723 -1688 -1689 -712
rect -1465 -1688 -1431 -712
rect 1431 -1688 1465 -712
rect 1689 -1688 1723 -712
rect -1611 -1772 -1543 -1738
rect -1396 -1772 -1342 -1738
rect -685 -1902 -605 -1822
rect -427 -1902 -347 -1822
rect 347 -1902 427 -1822
rect 605 -1902 685 -1822
rect 1342 -1772 1396 -1738
rect 1543 -1772 1611 -1738
rect -556 -2126 -476 -2046
rect 476 -2126 556 -2046
rect 2822 -4117 2922 -423
rect -2822 -4422 -2760 -4322
rect -2760 -4422 2760 -4322
rect 2760 -4422 2822 -4322
<< metal1 >>
rect -2928 4422 2928 4428
rect -2928 4322 -2822 4422
rect 2822 4322 2928 4422
rect -2928 4316 2928 4322
rect -2928 4117 -2816 4316
rect -2928 423 -2922 4117
rect -2822 3746 -2816 4117
rect -2216 4016 -2206 4316
rect 2206 4016 2216 4316
rect 2816 4117 2928 4316
rect 2816 3746 2822 4117
rect -2822 3654 -235 3746
rect -2822 2038 -2816 3654
rect -2345 3587 -2299 3654
rect -2345 3541 -2147 3587
rect -2345 3471 -2299 3541
rect -1829 3471 -1783 3654
rect -1313 3587 -1267 3654
rect -1313 3541 -1115 3587
rect -1313 3471 -1267 3541
rect -797 3471 -751 3654
rect -281 3471 -235 3654
rect 235 3654 2822 3746
rect 235 3500 281 3654
rect 751 3500 797 3654
rect 1267 3587 1313 3654
rect 1115 3541 1313 3587
rect 1267 3500 1313 3541
rect 1783 3500 1829 3654
rect 2299 3587 2345 3654
rect 2147 3541 2345 3587
rect 2299 3500 2345 3541
rect -2087 2459 -2041 2500
rect -2087 2367 -1889 2459
rect -2087 2162 -2041 2367
rect -1571 2254 -1525 2500
rect -1055 2459 -1009 2500
rect -1055 2367 -857 2459
rect -1571 2248 -1507 2254
rect -1571 2196 -1565 2248
rect -1513 2196 -1507 2248
rect -1571 2190 -1507 2196
rect -1055 2162 -1009 2367
rect -539 2346 -493 2500
rect -23 2459 23 2500
rect -175 2450 175 2459
rect -175 2389 -54 2450
rect 55 2389 175 2450
rect -175 2380 175 2389
rect 493 2346 539 2500
rect 1009 2459 1055 2500
rect 857 2367 1055 2459
rect -539 2340 -475 2346
rect -671 2288 -567 2294
rect -671 2196 -665 2288
rect -573 2196 -567 2288
rect -539 2288 -533 2340
rect -481 2288 -475 2340
rect -539 2282 -475 2288
rect -33 2340 31 2346
rect -33 2288 -27 2340
rect 25 2288 31 2340
rect -671 2190 -567 2196
rect -2087 2156 -2023 2162
rect -2087 2104 -2081 2156
rect -2029 2104 -2023 2156
rect -2087 2098 -2023 2104
rect -1064 2156 -1000 2162
rect -1064 2104 -1058 2156
rect -1006 2104 -1000 2156
rect -1064 2098 -1000 2104
rect -2822 2010 -1115 2038
rect -2822 1890 -2816 2010
rect -2556 1976 -1238 1982
rect -2556 1924 -2550 1976
rect -2498 1924 -1238 1976
rect -2556 1918 -1238 1924
rect -1302 1912 -1238 1918
rect -2822 1826 -1436 1890
rect -2822 423 -2816 1826
rect -1471 1787 -1436 1826
rect -1302 1860 -1296 1912
rect -1244 1860 -1238 1912
rect -1302 1854 -1238 1860
rect -1729 1781 -1436 1787
rect -1729 1747 -1611 1781
rect -1543 1747 -1436 1781
rect -1729 1741 -1436 1747
rect -1408 1781 -1330 1787
rect -1408 1747 -1396 1781
rect -1342 1747 -1330 1781
rect -1408 1741 -1330 1747
rect -1729 1688 -1683 1741
rect -1729 712 -1723 1688
rect -1689 712 -1683 1688
rect -1729 700 -1683 712
rect -1471 1700 -1436 1741
rect -1302 1700 -1267 1854
rect -1207 1741 -1115 2010
rect -975 2014 -901 2020
rect -975 1952 -969 2014
rect -907 1952 -901 2014
rect -975 1946 -901 1952
rect -797 2004 -733 2010
rect -797 1952 -791 2004
rect -739 1952 -733 2004
rect -797 1946 -733 1952
rect -290 2003 -226 2009
rect -290 1951 -284 2003
rect -232 1951 -226 2003
rect -797 1700 -751 1946
rect -290 1945 -226 1951
rect -33 2004 31 2288
rect 475 2340 539 2346
rect 475 2288 481 2340
rect 533 2288 539 2340
rect 475 2282 539 2288
rect 567 2288 671 2294
rect 567 2196 573 2288
rect 665 2196 671 2288
rect 567 2190 671 2196
rect 1009 2162 1055 2367
rect 1525 2254 1571 2500
rect 2041 2459 2087 2500
rect 1889 2367 2087 2459
rect 1507 2248 1571 2254
rect 1507 2196 1513 2248
rect 1565 2196 1571 2248
rect 1507 2190 1571 2196
rect 2041 2162 2087 2367
rect 1000 2156 1064 2162
rect 1000 2104 1006 2156
rect 1058 2104 1064 2156
rect 1000 2098 1064 2104
rect 2023 2156 2087 2162
rect 2023 2104 2029 2156
rect 2081 2104 2087 2156
rect 2023 2098 2087 2104
rect 2816 2038 2822 3654
rect 901 2014 975 2020
rect -33 1952 -27 2004
rect 25 1952 31 2004
rect -33 1945 31 1952
rect 226 2004 290 2010
rect 226 1952 232 2004
rect 284 1952 290 2004
rect 226 1946 290 1952
rect 733 2004 797 2010
rect 733 1952 739 2004
rect 791 1952 797 2004
rect 733 1946 797 1952
rect 901 1952 907 2014
rect 969 1952 975 2014
rect 901 1946 975 1952
rect 1115 2010 2822 2038
rect -1471 1688 -1425 1700
rect -1471 712 -1465 1688
rect -1431 712 -1425 1688
rect -281 1687 -235 1945
rect 235 1700 281 1946
rect 751 1700 797 1946
rect 1115 1741 1207 2010
rect 1238 1976 2551 1982
rect 1238 1924 2493 1976
rect 2545 1924 2551 1976
rect 1238 1918 2551 1924
rect 1238 1912 1302 1918
rect 1238 1860 1244 1912
rect 1296 1860 1302 1912
rect 2816 1890 2822 2010
rect 1238 1854 1302 1860
rect 1267 1700 1302 1854
rect 1436 1826 2822 1890
rect 1436 1787 1471 1826
rect 1330 1781 1408 1787
rect 1330 1747 1342 1781
rect 1396 1747 1408 1781
rect 1330 1741 1408 1747
rect 1436 1781 1729 1787
rect 1436 1747 1543 1781
rect 1611 1747 1729 1781
rect 1436 1741 1729 1747
rect 1436 1700 1471 1741
rect 1425 1688 1471 1700
rect -1471 700 -1425 712
rect 1425 712 1431 1688
rect 1465 712 1471 1688
rect 1425 700 1471 712
rect 1683 1688 1729 1741
rect 1683 712 1689 1688
rect 1723 712 1729 1688
rect 1683 700 1729 712
rect -1623 653 -1531 659
rect -1623 619 -1611 653
rect -1543 619 -1531 653
rect -1623 613 -1531 619
rect -1408 653 -1330 659
rect -1408 619 -1396 653
rect -1342 619 -1330 653
rect -1408 613 -1330 619
rect -1274 573 -1200 579
rect -1274 511 -1268 573
rect -1206 511 -1200 573
rect -1274 505 -1200 511
rect -1055 546 -1009 700
rect -1055 540 -991 546
rect -1055 488 -1049 540
rect -997 488 -991 540
rect -1055 482 -991 488
rect -2928 224 -2816 423
rect -539 362 -493 700
rect -23 546 23 700
rect -32 540 32 546
rect -32 488 -26 540
rect 26 488 32 540
rect -32 482 32 488
rect 493 362 539 700
rect 1009 546 1055 700
rect 1330 653 1408 659
rect 1330 619 1342 653
rect 1396 619 1408 653
rect 1330 613 1408 619
rect 1531 653 1623 659
rect 1531 619 1543 653
rect 1611 619 1623 653
rect 1531 613 1623 619
rect 991 540 1055 546
rect 991 488 997 540
rect 1049 488 1055 540
rect 1190 573 1264 579
rect 1190 511 1196 573
rect 1258 511 1264 573
rect 1190 505 1264 511
rect 991 482 1055 488
rect 2816 423 2822 1826
rect 2922 423 2928 4117
rect -2392 356 -475 362
rect -2392 304 -2386 356
rect -2334 304 -533 356
rect -481 304 -475 356
rect -2392 298 -475 304
rect 475 356 2391 362
rect 475 304 481 356
rect 533 304 2333 356
rect 2385 304 2391 356
rect 475 298 2391 304
rect 2816 224 2928 423
rect -2928 218 2928 224
rect -2928 118 -2822 218
rect 2822 118 2928 218
rect -2928 112 2928 118
rect -2928 -118 2928 -112
rect -2928 -218 -2822 -118
rect 2822 -218 2928 -118
rect -2928 -224 2928 -218
rect -2928 -252 -2816 -224
rect 2816 -252 2928 -224
rect -2928 -316 2928 -252
rect -2928 -423 -2816 -316
rect -2556 -360 -1672 -354
rect -2556 -412 -2550 -360
rect -2498 -412 -1730 -360
rect -1678 -412 -1672 -360
rect -2556 -418 -1672 -412
rect -2928 -4117 -2922 -423
rect -2822 -2166 -2816 -423
rect -1471 -622 -1436 -316
rect -1302 -360 -1238 -354
rect -1302 -412 -1296 -360
rect -1244 -412 -1238 -360
rect -1302 -418 -1238 -412
rect -1729 -628 -1436 -622
rect -1729 -662 -1611 -628
rect -1543 -662 -1436 -628
rect -1729 -668 -1436 -662
rect -1408 -628 -1330 -622
rect -1408 -662 -1396 -628
rect -1342 -662 -1330 -628
rect -1408 -668 -1330 -662
rect -1729 -712 -1683 -668
rect -1729 -1688 -1723 -712
rect -1689 -1688 -1683 -712
rect -1729 -1700 -1683 -1688
rect -1471 -700 -1436 -668
rect -1302 -700 -1267 -418
rect -1207 -668 -1115 -316
rect -797 -700 -751 -316
rect -281 -700 -235 -316
rect -199 -360 207 -354
rect -199 -412 -193 -360
rect -141 -412 149 -360
rect 201 -412 207 -360
rect -199 -418 207 -412
rect -53 -452 51 -446
rect -53 -544 -47 -452
rect 45 -544 51 -452
rect -53 -550 51 -544
rect 235 -700 281 -316
rect 751 -700 797 -316
rect 1115 -668 1207 -316
rect 1238 -360 1302 -354
rect 1238 -412 1244 -360
rect 1296 -412 1302 -360
rect 1238 -418 1302 -412
rect 1267 -700 1302 -418
rect 1436 -622 1471 -316
rect 1671 -360 2551 -354
rect 1671 -412 1677 -360
rect 1729 -412 2493 -360
rect 2545 -412 2551 -360
rect 1671 -418 2551 -412
rect 2816 -423 2928 -316
rect 1330 -628 1408 -622
rect 1330 -662 1342 -628
rect 1396 -662 1408 -628
rect 1330 -668 1408 -662
rect 1436 -628 1729 -622
rect 1436 -662 1543 -628
rect 1611 -662 1729 -628
rect 1436 -668 1729 -662
rect 1436 -700 1471 -668
rect -1471 -712 -1425 -700
rect -1471 -1688 -1465 -712
rect -1431 -1688 -1425 -712
rect -1471 -1700 -1425 -1688
rect 1425 -712 1471 -700
rect 1425 -1688 1431 -712
rect 1465 -1688 1471 -712
rect 1425 -1700 1471 -1688
rect 1683 -712 1729 -668
rect 1683 -1688 1689 -712
rect 1723 -1688 1729 -712
rect 1683 -1700 1729 -1688
rect -1623 -1738 -1531 -1732
rect -1623 -1772 -1611 -1738
rect -1543 -1772 -1531 -1738
rect -1623 -1778 -1531 -1772
rect -1408 -1738 -1330 -1732
rect -1408 -1772 -1396 -1738
rect -1342 -1772 -1330 -1738
rect -1408 -1778 -1330 -1772
rect -2556 -1856 -1836 -1850
rect -2556 -1908 -2550 -1856
rect -2498 -1908 -1894 -1856
rect -1842 -1908 -1836 -1856
rect -2556 -1914 -1836 -1908
rect -1055 -2034 -1009 -1700
rect -697 -1816 -593 -1810
rect -697 -1908 -691 -1816
rect -599 -1908 -593 -1816
rect -697 -1914 -593 -1908
rect -539 -1942 -493 -1700
rect -439 -1816 -335 -1810
rect -439 -1908 -433 -1816
rect -341 -1908 -335 -1816
rect -439 -1914 -335 -1908
rect -539 -1948 -475 -1942
rect -539 -2000 -533 -1948
rect -481 -2000 -475 -1948
rect -539 -2006 -475 -2000
rect -23 -2034 23 -1700
rect 335 -1816 439 -1810
rect 335 -1908 341 -1816
rect 433 -1908 439 -1816
rect 335 -1914 439 -1908
rect 493 -1942 539 -1700
rect 593 -1816 697 -1810
rect 593 -1908 599 -1816
rect 691 -1908 697 -1816
rect 593 -1914 697 -1908
rect 475 -1948 539 -1942
rect 475 -2000 481 -1948
rect 533 -2000 539 -1948
rect 475 -2006 539 -2000
rect 1009 -2034 1055 -1700
rect 1330 -1738 1408 -1732
rect 1330 -1772 1342 -1738
rect 1396 -1772 1408 -1738
rect 1330 -1778 1408 -1772
rect 1531 -1738 1623 -1732
rect 1531 -1772 1543 -1738
rect 1611 -1772 1623 -1738
rect 1531 -1778 1623 -1772
rect 1835 -1856 2555 -1850
rect 1835 -1908 1841 -1856
rect 1893 -1908 2497 -1856
rect 2549 -1908 2555 -1856
rect 1835 -1914 2555 -1908
rect -1055 -2040 -991 -2034
rect -1055 -2092 -1049 -2040
rect -997 -2092 -991 -2040
rect -1055 -2098 -991 -2092
rect -568 -2040 -464 -2034
rect -568 -2132 -562 -2040
rect -470 -2132 -464 -2040
rect -32 -2040 32 -2034
rect -32 -2092 -26 -2040
rect 26 -2092 32 -2040
rect -32 -2098 32 -2092
rect 464 -2040 568 -2034
rect -568 -2138 -464 -2132
rect 464 -2132 470 -2040
rect 562 -2132 568 -2040
rect 991 -2040 1055 -2034
rect 991 -2092 997 -2040
rect 1049 -2092 1055 -2040
rect 991 -2098 1055 -2092
rect 464 -2138 568 -2132
rect 2816 -2166 2822 -423
rect -2822 -2230 2822 -2166
rect -2822 -4117 -2816 -2230
rect -2239 -2428 -2147 -2230
rect -2096 -2316 -2032 -2310
rect -2096 -2368 -2090 -2316
rect -2038 -2368 -2032 -2316
rect -2096 -2374 -2032 -2368
rect -2345 -2468 -2147 -2428
rect -2345 -2500 -2299 -2468
rect -2087 -2500 -2041 -2374
rect -1829 -2500 -1783 -2230
rect -1723 -2316 -1631 -2310
rect -1723 -2368 -1717 -2316
rect -1637 -2368 -1631 -2316
rect -1723 -2468 -1631 -2368
rect -1465 -2316 -1373 -2310
rect -1465 -2368 -1459 -2316
rect -1379 -2368 -1373 -2316
rect -1465 -2468 -1373 -2368
rect -1313 -2500 -1267 -2230
rect -1064 -2316 -1000 -2310
rect -1064 -2368 -1058 -2316
rect -1006 -2368 -1000 -2316
rect -1064 -2374 -1000 -2368
rect -1055 -2500 -1009 -2374
rect -949 -2468 -857 -2230
rect -539 -2500 -493 -2230
rect -433 -2316 -341 -2310
rect -433 -2368 -427 -2316
rect -347 -2368 -341 -2316
rect -433 -2412 -341 -2368
rect -290 -2316 -226 -2310
rect -290 -2368 -284 -2316
rect -232 -2368 -226 -2316
rect -290 -2374 -226 -2368
rect -175 -2316 -83 -2310
rect -175 -2368 -169 -2316
rect -89 -2368 -83 -2316
rect -281 -2412 -235 -2374
rect -175 -2412 -83 -2368
rect -433 -2468 -83 -2412
rect -281 -2500 -235 -2468
rect -23 -2500 23 -2230
rect 493 -2500 539 -2230
rect 599 -2316 691 -2310
rect 599 -2368 605 -2316
rect 685 -2368 691 -2316
rect 599 -2412 691 -2368
rect 742 -2316 806 -2310
rect 742 -2368 748 -2316
rect 800 -2368 806 -2316
rect 742 -2374 806 -2368
rect 751 -2412 797 -2374
rect 599 -2468 797 -2412
rect 857 -2468 949 -2230
rect 1000 -2316 1064 -2310
rect 1000 -2368 1006 -2316
rect 1058 -2368 1064 -2316
rect 1000 -2374 1064 -2368
rect 751 -2500 797 -2468
rect 1009 -2500 1055 -2374
rect 1267 -2500 1313 -2230
rect 1373 -2316 1465 -2310
rect 1373 -2368 1379 -2316
rect 1459 -2368 1465 -2316
rect 1373 -2468 1465 -2368
rect 1631 -2316 1723 -2310
rect 1631 -2368 1637 -2316
rect 1717 -2368 1723 -2316
rect 1631 -2468 1723 -2368
rect 1783 -2500 1829 -2230
rect 2032 -2316 2096 -2310
rect 2032 -2368 2038 -2316
rect 2090 -2368 2096 -2316
rect 2032 -2374 2096 -2368
rect 2041 -2500 2087 -2374
rect 2147 -2428 2239 -2230
rect 2147 -2468 2345 -2428
rect 2299 -2500 2345 -2468
rect -1981 -3632 -1889 -3532
rect -1571 -3626 -1525 -3500
rect -797 -3532 -751 -3500
rect 235 -3532 281 -3500
rect -1981 -3684 -1975 -3632
rect -1895 -3684 -1889 -3632
rect -1981 -3690 -1889 -3684
rect -1580 -3632 -1516 -3626
rect -1580 -3684 -1574 -3632
rect -1522 -3684 -1516 -3632
rect -1580 -3690 -1516 -3684
rect -1207 -3632 -1115 -3532
rect -797 -3588 -599 -3532
rect -797 -3626 -751 -3588
rect -1207 -3684 -1201 -3632
rect -1121 -3684 -1115 -3632
rect -1207 -3690 -1115 -3684
rect -806 -3632 -742 -3626
rect -806 -3684 -800 -3632
rect -748 -3684 -742 -3632
rect -806 -3690 -742 -3684
rect -691 -3632 -599 -3588
rect -691 -3684 -685 -3632
rect -605 -3684 -599 -3632
rect -691 -3690 -599 -3684
rect 83 -3589 433 -3532
rect 83 -3632 175 -3589
rect 235 -3626 281 -3589
rect 83 -3684 89 -3632
rect 169 -3684 175 -3632
rect 83 -3690 175 -3684
rect 226 -3632 290 -3626
rect 226 -3684 232 -3632
rect 284 -3684 290 -3632
rect 226 -3690 290 -3684
rect 341 -3632 433 -3589
rect 341 -3684 347 -3632
rect 427 -3684 433 -3632
rect 341 -3690 433 -3684
rect 1115 -3632 1207 -3532
rect 1525 -3626 1571 -3500
rect 1115 -3684 1121 -3632
rect 1201 -3684 1207 -3632
rect 1115 -3690 1207 -3684
rect 1516 -3632 1580 -3626
rect 1516 -3684 1522 -3632
rect 1574 -3684 1580 -3632
rect 1516 -3690 1580 -3684
rect 1889 -3632 1981 -3532
rect 1889 -3684 1895 -3632
rect 1975 -3684 1981 -3632
rect 1889 -3690 1981 -3684
rect -2928 -4316 -2816 -4117
rect -2216 -4316 -2206 -4016
rect 2206 -4316 2216 -4016
rect 2816 -4117 2822 -2230
rect 2922 -4117 2928 -423
rect 2816 -4316 2928 -4117
rect -2928 -4322 2928 -4316
rect -2928 -4422 -2822 -4322
rect 2822 -4422 2928 -4322
rect -2928 -4428 2928 -4422
<< via1 >>
rect -2816 4016 -2216 4316
rect 2216 4016 2816 4316
rect -1565 2196 -1513 2248
rect -54 2389 55 2450
rect -665 2282 -573 2288
rect -665 2202 -659 2282
rect -659 2202 -579 2282
rect -579 2202 -573 2282
rect -665 2196 -573 2202
rect -533 2288 -481 2340
rect -27 2288 25 2340
rect -2081 2104 -2029 2156
rect -1058 2104 -1006 2156
rect -2550 1924 -2498 1976
rect -1296 1860 -1244 1912
rect -969 2008 -907 2014
rect -969 1958 -963 2008
rect -963 1958 -913 2008
rect -913 1958 -907 2008
rect -969 1952 -907 1958
rect -791 1952 -739 2004
rect -284 1951 -232 2003
rect 481 2288 533 2340
rect 573 2282 665 2288
rect 573 2202 579 2282
rect 579 2202 659 2282
rect 659 2202 665 2282
rect 573 2196 665 2202
rect 1513 2196 1565 2248
rect 1006 2104 1058 2156
rect 2029 2104 2081 2156
rect -27 1952 25 2004
rect 232 1952 284 2004
rect 739 1952 791 2004
rect 907 2008 969 2014
rect 907 1958 913 2008
rect 913 1958 963 2008
rect 963 1958 969 2008
rect 907 1952 969 1958
rect 2493 1924 2545 1976
rect 1244 1860 1296 1912
rect -1268 567 -1206 573
rect -1268 517 -1262 567
rect -1262 517 -1212 567
rect -1212 517 -1206 567
rect -1268 511 -1206 517
rect -1049 488 -997 540
rect -26 488 26 540
rect 997 488 1049 540
rect 1196 567 1258 573
rect 1196 517 1202 567
rect 1202 517 1252 567
rect 1252 517 1258 567
rect 1196 511 1258 517
rect -2386 304 -2334 356
rect -533 304 -481 356
rect 481 304 533 356
rect 2333 304 2385 356
rect -2550 -412 -2498 -360
rect -1730 -412 -1678 -360
rect -1296 -412 -1244 -360
rect -193 -412 -141 -360
rect 149 -412 201 -360
rect -47 -458 45 -452
rect -47 -538 -41 -458
rect -41 -538 39 -458
rect 39 -538 45 -458
rect -47 -544 45 -538
rect 1244 -412 1296 -360
rect 1677 -412 1729 -360
rect 2493 -412 2545 -360
rect -2550 -1908 -2498 -1856
rect -1894 -1908 -1842 -1856
rect -691 -1822 -599 -1816
rect -691 -1902 -685 -1822
rect -685 -1902 -605 -1822
rect -605 -1902 -599 -1822
rect -691 -1908 -599 -1902
rect -433 -1822 -341 -1816
rect -433 -1902 -427 -1822
rect -427 -1902 -347 -1822
rect -347 -1902 -341 -1822
rect -433 -1908 -341 -1902
rect -533 -2000 -481 -1948
rect 341 -1822 433 -1816
rect 341 -1902 347 -1822
rect 347 -1902 427 -1822
rect 427 -1902 433 -1822
rect 341 -1908 433 -1902
rect 599 -1822 691 -1816
rect 599 -1902 605 -1822
rect 605 -1902 685 -1822
rect 685 -1902 691 -1822
rect 599 -1908 691 -1902
rect 481 -2000 533 -1948
rect 1841 -1908 1893 -1856
rect 2497 -1908 2549 -1856
rect -1049 -2092 -997 -2040
rect -562 -2046 -470 -2040
rect -562 -2126 -556 -2046
rect -556 -2126 -476 -2046
rect -476 -2126 -470 -2046
rect -562 -2132 -470 -2126
rect -26 -2092 26 -2040
rect 470 -2046 562 -2040
rect 470 -2126 476 -2046
rect 476 -2126 556 -2046
rect 556 -2126 562 -2046
rect 470 -2132 562 -2126
rect 997 -2092 1049 -2040
rect -2090 -2368 -2038 -2316
rect -1717 -2368 -1637 -2316
rect -1459 -2368 -1379 -2316
rect -1058 -2368 -1006 -2316
rect -427 -2368 -347 -2316
rect -284 -2368 -232 -2316
rect -169 -2368 -89 -2316
rect 605 -2368 685 -2316
rect 748 -2368 800 -2316
rect 1006 -2368 1058 -2316
rect 1379 -2368 1459 -2316
rect 1637 -2368 1717 -2316
rect 2038 -2368 2090 -2316
rect -1975 -3684 -1895 -3632
rect -1574 -3684 -1522 -3632
rect -1201 -3684 -1121 -3632
rect -800 -3684 -748 -3632
rect -685 -3684 -605 -3632
rect 89 -3684 169 -3632
rect 232 -3684 284 -3632
rect 347 -3684 427 -3632
rect 1121 -3684 1201 -3632
rect 1522 -3684 1574 -3632
rect 1895 -3684 1975 -3632
rect -2816 -4316 -2216 -4016
rect 2216 -4316 2816 -4016
<< metal2 >>
rect -2816 4316 -2216 4326
rect -2816 4006 -2216 4016
rect 2216 4316 2816 4326
rect 2216 4006 2816 4016
rect -63 2450 63 2459
rect -63 2389 -54 2450
rect 55 2389 63 2450
rect -63 2380 63 2389
rect -539 2340 539 2346
rect -671 2288 -567 2294
rect -671 2254 -665 2288
rect -2228 2248 -665 2254
rect -2228 2196 -1565 2248
rect -1513 2196 -665 2248
rect -573 2254 -567 2288
rect -539 2288 -533 2340
rect -481 2288 -27 2340
rect 25 2288 481 2340
rect 533 2288 539 2340
rect -539 2282 539 2288
rect 567 2288 671 2294
rect 567 2254 573 2288
rect -573 2196 573 2254
rect 665 2254 671 2288
rect 665 2248 2227 2254
rect 665 2196 1513 2248
rect 1565 2196 2227 2248
rect -2228 2190 2227 2196
rect -2556 1976 -2492 1982
rect -2556 1924 -2550 1976
rect -2498 1924 -2492 1976
rect -2556 -360 -2492 1924
rect -2556 -412 -2550 -360
rect -2498 -412 -2492 -360
rect -2556 -418 -2492 -412
rect -2392 356 -2328 362
rect -2392 304 -2386 356
rect -2334 304 -2328 356
rect -2556 -1856 -2492 -1850
rect -2556 -1908 -2550 -1856
rect -2498 -1908 -2492 -1856
rect -2556 -3718 -2492 -1908
rect -2392 -2218 -2328 304
rect -2228 -2034 -2164 2190
rect -2087 2156 2087 2162
rect -2087 2104 -2081 2156
rect -2029 2104 -1058 2156
rect -1006 2104 1006 2156
rect 1058 2104 2029 2156
rect 2081 2104 2087 2156
rect -2087 2098 2087 2104
rect -1576 2070 -1512 2098
rect -2064 2006 -1512 2070
rect 1512 2070 1576 2098
rect -975 2014 -901 2020
rect -2064 -1942 -2000 2006
rect -975 1952 -969 2014
rect -907 1952 -901 2014
rect 901 2014 975 2020
rect -975 1946 -901 1952
rect -797 2004 797 2010
rect -797 1952 -791 2004
rect -739 2003 -27 2004
rect -739 1952 -284 2003
rect -797 1951 -284 1952
rect -232 1952 -27 2003
rect 25 1952 232 2004
rect 284 1952 739 2004
rect 791 1952 797 2004
rect -232 1951 797 1952
rect -797 1946 797 1951
rect 901 1952 907 2014
rect 969 1952 975 2014
rect 1512 2006 2063 2070
rect 901 1946 975 1952
rect -1302 1912 1302 1918
rect -1302 1860 -1296 1912
rect -1244 1860 1244 1912
rect 1296 1860 1302 1912
rect -1302 1854 1302 1860
rect -1274 573 -1200 579
rect -1274 511 -1268 573
rect -1206 511 -1200 573
rect 1190 573 1264 579
rect -1274 505 -1200 511
rect -1055 540 1055 546
rect -1055 488 -1049 540
rect -997 488 -26 540
rect 26 488 997 540
rect 1049 488 1055 540
rect 1190 511 1196 573
rect 1258 511 1264 573
rect 1190 505 1264 511
rect -1055 482 1055 488
rect -32 454 32 482
rect -1900 390 1899 454
rect -1900 -1850 -1836 390
rect -539 356 539 362
rect -539 304 -533 356
rect -481 304 481 356
rect 533 304 539 356
rect -539 298 539 304
rect -1736 -360 -135 -354
rect -1736 -412 -1730 -360
rect -1678 -412 -1296 -360
rect -1244 -412 -193 -360
rect -141 -412 -135 -360
rect -1736 -418 -135 -412
rect -33 -446 31 298
rect 143 -360 1735 -354
rect 143 -412 149 -360
rect 201 -412 1244 -360
rect 1296 -412 1677 -360
rect 1729 -412 1735 -360
rect 143 -418 1735 -412
rect -53 -452 51 -446
rect -53 -544 -47 -452
rect 45 -544 51 -452
rect -53 -550 51 -544
rect -697 -1816 -593 -1810
rect -697 -1850 -691 -1816
rect -1900 -1856 -691 -1850
rect -1900 -1908 -1894 -1856
rect -1842 -1908 -691 -1856
rect -599 -1850 -593 -1816
rect -439 -1816 -335 -1810
rect -439 -1850 -433 -1816
rect -599 -1908 -433 -1850
rect -341 -1908 -335 -1816
rect -1900 -1914 -335 -1908
rect 335 -1816 439 -1810
rect 335 -1908 341 -1816
rect 433 -1850 439 -1816
rect 593 -1816 697 -1810
rect 593 -1850 599 -1816
rect 433 -1908 599 -1850
rect 691 -1850 697 -1816
rect 1835 -1850 1899 390
rect 691 -1856 1899 -1850
rect 691 -1908 1841 -1856
rect 1893 -1908 1899 -1856
rect 335 -1914 1899 -1908
rect 1999 -1942 2063 2006
rect -2064 -1948 2063 -1942
rect -2064 -2000 -533 -1948
rect -481 -2000 481 -1948
rect 533 -2000 2063 -1948
rect -2064 -2006 2063 -2000
rect 2163 -2034 2227 2190
rect 2487 1976 2551 1982
rect 2487 1924 2493 1976
rect 2545 1924 2551 1976
rect 2487 819 2551 1924
rect 2482 810 2556 819
rect 2482 754 2491 810
rect 2547 754 2556 810
rect 2482 745 2556 754
rect -2228 -2040 2227 -2034
rect -2228 -2092 -1049 -2040
rect -997 -2092 -562 -2040
rect -2228 -2098 -562 -2092
rect -568 -2132 -562 -2098
rect -470 -2092 -26 -2040
rect 26 -2092 470 -2040
rect -470 -2098 470 -2092
rect -470 -2132 -464 -2098
rect -568 -2138 -464 -2132
rect 464 -2132 470 -2098
rect 562 -2092 997 -2040
rect 1049 -2092 2227 -2040
rect 562 -2098 2227 -2092
rect 2327 356 2391 362
rect 2327 304 2333 356
rect 2385 304 2391 356
rect 562 -2132 568 -2098
rect 464 -2138 568 -2132
rect 2327 -2218 2391 304
rect 2487 -360 2551 745
rect 2487 -412 2493 -360
rect 2545 -412 2551 -360
rect 2487 -418 2551 -412
rect -2392 -2282 2391 -2218
rect 2491 -1856 2555 -1850
rect 2491 -1908 2497 -1856
rect 2549 -1908 2555 -1856
rect 2491 -1933 2555 -1908
rect -32 -2310 32 -2282
rect -2096 -2316 2096 -2310
rect -2096 -2368 -2090 -2316
rect -2038 -2368 -1717 -2316
rect -1637 -2368 -1459 -2316
rect -1379 -2368 -1058 -2316
rect -1006 -2368 -427 -2316
rect -347 -2368 -284 -2316
rect -232 -2368 -169 -2316
rect -89 -2368 605 -2316
rect 685 -2368 748 -2316
rect 800 -2368 1006 -2316
rect 1058 -2368 1379 -2316
rect 1459 -2368 1637 -2316
rect 1717 -2368 2038 -2316
rect 2090 -2368 2096 -2316
rect -2096 -2374 2096 -2368
rect -1981 -3632 1981 -3626
rect -1981 -3684 -1975 -3632
rect -1895 -3684 -1574 -3632
rect -1522 -3684 -1201 -3632
rect -1121 -3684 -800 -3632
rect -748 -3684 -685 -3632
rect -605 -3684 89 -3632
rect 169 -3684 232 -3632
rect 284 -3684 347 -3632
rect 427 -3684 1121 -3632
rect 1201 -3684 1522 -3632
rect 1574 -3684 1895 -3632
rect 1975 -3684 1981 -3632
rect -1981 -3690 1981 -3684
rect -32 -3718 32 -3690
rect 2491 -3718 2556 -1933
rect -2556 -3782 2556 -3718
rect -2816 -4016 -2216 -4006
rect -2816 -4326 -2216 -4316
rect 2216 -4016 2816 -4006
rect 2216 -4326 2816 -4316
<< via2 >>
rect -2816 4016 -2216 4316
rect 2216 4016 2816 4316
rect -54 2389 55 2450
rect -966 1955 -910 2011
rect 910 1955 966 2011
rect -1265 514 -1209 570
rect 1199 514 1255 570
rect 2491 754 2547 810
rect -2816 -4316 -2216 -4016
rect 2216 -4316 2816 -4016
<< metal3 >>
rect -2826 4316 -2206 4321
rect -2826 4016 -2816 4316
rect -2216 4016 -2206 4316
rect -2826 4011 -2206 4016
rect 2206 4316 2826 4321
rect 2206 4016 2216 4316
rect 2816 4016 2826 4316
rect 2206 4011 2826 4016
rect -63 2450 63 2459
rect -63 2389 -54 2450
rect 55 2389 63 2450
rect -63 2380 63 2389
rect -2595 2320 63 2380
rect -2595 2153 50 2213
rect -50 2093 50 2153
rect -988 2033 988 2093
rect -988 2011 -888 2033
rect -988 1955 -966 2011
rect -910 1955 -888 2011
rect -988 1933 -888 1955
rect 888 2011 988 2033
rect 888 1955 910 2011
rect 966 1955 988 2011
rect 888 1933 988 1955
rect 2469 812 2569 832
rect 2469 810 2737 812
rect 2469 754 2491 810
rect 2547 754 2737 810
rect 2469 752 2737 754
rect 2469 732 2569 752
rect -1287 570 -1187 592
rect -1287 514 -1265 570
rect -1209 514 -1187 570
rect -1287 492 -1187 514
rect 1177 570 1277 592
rect 1177 514 1199 570
rect 1255 514 1277 570
rect 1177 492 1277 514
rect -1287 432 1277 492
rect -55 372 45 432
rect -2621 312 45 372
rect -2826 -4016 -2206 -4011
rect -2826 -4316 -2816 -4016
rect -2216 -4316 -2206 -4016
rect -2826 -4321 -2206 -4316
rect 2206 -4016 2826 -4011
rect 2206 -4316 2216 -4016
rect 2816 -4316 2826 -4016
rect 2206 -4321 2826 -4316
<< via3 >>
rect -2816 4016 -2216 4316
rect 2216 4016 2816 4316
rect -2816 -4316 -2216 -4016
rect 2216 -4316 2816 -4016
<< metal4 >>
rect -3000 4316 3000 4500
rect -3000 4016 -2816 4316
rect -2216 4016 2216 4316
rect 2816 4016 3000 4316
rect -3000 3700 3000 4016
rect -3000 -4016 3000 -3700
rect -3000 -4316 -2816 -4016
rect -2216 -4316 2216 -4016
rect 2816 -4316 3000 -4016
rect -3000 -4500 3000 -4316
use sky130_fd_pr__nfet_g5v0d10v5_V2YKKA  xm1 ../comparator
timestamp 1621838304
transform 1 0 0 0 1 -1200
box -1319 -588 1319 588
use sky130_fd_pr__nfet_g5v0d10v5_7QEKRB  xm2 ../comparator
timestamp 1621838304
transform 1 0 0 0 1 -3000
box -2351 -588 2351 588
use sky130_fd_pr__pfet_g5v0d10v5_QRGZLW  xm3 ../comparator
timestamp 1621838304
transform 1 0 0 0 1 1200
box -1385 -600 1385 600
use sky130_fd_pr__pfet_g5v0d10v5_QM5ZLW  xm4 ./../comparator
timestamp 1621838304
transform 1 0 0 0 1 3000
box -2417 -600 2417 600
<< labels >>
flabel metal4 -3000 3700 -3000 4500 3 FreeSans 480 0 0 0 vdd
port 2 e
flabel metal3 -2595 2153 -2595 2213 1 FreeSans 280 0 0 0 vinp
port 4 n
flabel metal3 -2621 312 -2621 372 1 FreeSans 280 0 0 0 vinm
port 3 n
flabel metal3 2737 752 2737 812 1 FreeSans 280 0 0 0 vout
port 5 n
flabel metal4 -3000 -4500 -2999 -3700 3 FreeSans 240 0 0 0 vss
port 6 e
flabel metal3 -2595 2320 -2595 2380 1 FreeSans 240 0 0 0 ibias
port 1 n
<< properties >>
string FIXED_BBOX -2872 -4372 2872 -168
<< end >>
