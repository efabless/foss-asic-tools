magic
tech sky130A
magscale 1 2
timestamp 1624430562
<< metal1 >>
rect 483489 547727 483495 547730
rect 447081 547681 483495 547727
rect 447081 547118 447127 547681
rect 483489 547678 483495 547681
rect 483547 547678 483553 547730
rect 446849 547072 447127 547118
rect 482910 547044 482916 547047
rect 446849 546998 482916 547044
rect 438114 546992 438204 546998
rect 482910 546995 482916 546998
rect 482968 546995 482974 547047
rect 438204 546970 441008 546992
rect 438204 546924 441423 546970
rect 438204 546902 441008 546924
rect 438114 546896 438204 546902
rect 447419 544531 447471 544537
rect 446849 544482 447419 544528
rect 438590 544387 438596 544475
rect 438684 544454 441067 544475
rect 447419 544473 447471 544479
rect 438684 544408 441423 544454
rect 446849 544408 447216 544454
rect 438684 544387 441067 544408
rect 447170 544400 447216 544408
rect 447245 544400 447251 544403
rect 447170 544354 447251 544400
rect 447245 544351 447251 544354
rect 447303 544351 447309 544403
rect 439085 541900 439202 541906
rect 439202 541818 441423 541864
rect 439085 541777 439202 541783
rect 439823 541438 439904 541444
rect 439904 541374 441423 541420
rect 439823 541351 439904 541357
rect 8448 537274 8454 541333
rect 12513 537274 16884 541333
rect 439548 541223 439644 541229
rect 439644 541152 441446 541198
rect 439548 541121 439644 541127
rect 440090 540980 440096 541065
rect 440181 541050 440336 541065
rect 440181 541004 441446 541050
rect 440181 540980 440336 541004
rect 437454 540830 437549 540836
rect 437549 540805 441073 540830
rect 437549 540759 441239 540805
rect 437549 540735 441073 540759
rect 437454 540729 437549 540735
rect 441193 540680 441239 540759
rect 441193 540634 441423 540680
rect 430931 540609 430983 540615
rect 430983 540560 441423 540606
rect 430931 540551 430983 540557
rect 441199 540486 441423 540532
rect 430631 540423 430683 540429
rect 441199 540420 441245 540486
rect 430683 540374 441245 540420
rect 430631 540365 430683 540371
rect 437016 539888 437103 539894
rect 437103 539801 440907 539888
rect 437016 539795 437103 539801
rect 440840 539749 440886 539801
rect 440840 539703 441142 539749
rect 441096 539644 441142 539703
rect 433176 539600 433281 539606
rect 433281 539570 440459 539600
rect 441096 539598 441423 539644
rect 447065 539570 447176 539576
rect 433281 539524 441423 539570
rect 446849 539524 447176 539570
rect 433281 539495 440459 539524
rect 447065 539516 447176 539524
rect 447236 539516 447242 539576
rect 433176 539489 433281 539495
rect 440914 539450 441423 539496
rect 440543 539052 440630 539058
rect 440914 539052 440960 539450
rect 440630 538965 440981 539052
rect 440543 538959 440630 538965
rect 1489 214412 7176 346469
rect 1489 210759 2293 214412
rect 5870 210759 7176 214412
rect 1489 18800 7176 210759
rect 12825 18800 16884 537274
<< via1 >>
rect 483495 547678 483547 547730
rect 482916 546995 482968 547047
rect 438114 546902 438204 546992
rect 447419 544479 447471 544531
rect 438596 544387 438684 544475
rect 447251 544351 447303 544403
rect 439085 541783 439202 541900
rect 439823 541357 439904 541438
rect 8454 537274 12513 541333
rect 439548 541127 439644 541223
rect 440096 540980 440181 541065
rect 437454 540735 437549 540830
rect 430931 540557 430983 540609
rect 430631 540371 430683 540423
rect 437016 539801 437103 539888
rect 433176 539495 433281 539600
rect 447176 539516 447236 539576
rect 440543 538965 440630 539052
rect 2293 210759 5870 214412
<< metal2 >>
rect 170894 701000 173094 701100
rect 170894 700500 170994 701000
rect 172994 700500 173094 701000
rect 170894 698400 173094 700500
rect 222594 701000 224794 701100
rect 222594 700500 222694 701000
rect 224694 700500 224794 701000
rect 222594 698400 224794 700500
rect 324294 701000 326494 701100
rect 324294 700500 324394 701000
rect 326394 700500 326494 701000
rect 324294 698400 326494 700500
rect 170894 587710 378401 698400
rect 576957 586033 577069 586038
rect 576953 585931 576962 586033
rect 577064 585931 577073 586033
rect 446924 555365 446970 555867
rect 447288 555622 447334 555830
rect 447288 555576 447468 555622
rect 446924 555319 447300 555365
rect 446174 549540 446874 549600
rect 446174 548061 446236 549540
rect 446814 548061 446874 549540
rect 438108 546902 438114 546992
rect 438204 546902 438210 546992
rect 446174 546957 446874 548061
rect 430909 545126 430987 545130
rect 430904 545121 430992 545126
rect 430904 545043 430909 545121
rect 430987 545043 430992 545121
rect 430904 544989 430992 545043
rect 430628 544334 430684 544341
rect 430626 544332 430686 544334
rect 430626 544276 430628 544332
rect 430684 544276 430686 544332
rect 430626 544234 430686 544276
rect 23814 543501 23823 543701
rect 24023 543501 24032 543701
rect 8454 541333 12513 541339
rect 5902 537274 5911 541333
rect 8454 537268 12513 537274
rect 11300 523331 11560 523336
rect 11296 523081 11305 523331
rect 11555 523081 11564 523331
rect 6816 509177 6825 509271
rect 6919 509177 6928 509271
rect 6825 481874 6919 509177
rect 6821 481790 6830 481874
rect 6914 481790 6923 481874
rect 6825 481785 6919 481790
rect 5291 480673 5378 480678
rect 5287 480596 5296 480673
rect 5373 480596 5382 480673
rect 3071 479741 3158 479746
rect 3067 479664 3076 479741
rect 3153 479664 3162 479741
rect 3071 422824 3158 479664
rect 5291 466063 5378 480596
rect 5282 465976 5291 466063
rect 5378 465976 5387 466063
rect 3062 422737 3071 422824
rect 3158 422737 3167 422824
rect 11300 382087 11560 523081
rect 15780 510027 15880 510032
rect 15776 509937 15785 510027
rect 15875 509937 15884 510027
rect 13406 507910 13606 507915
rect 13402 507720 13411 507910
rect 13601 507720 13610 507910
rect 11300 381818 11560 381827
rect 13406 350570 13606 507720
rect 9843 350370 13606 350570
rect 9843 345692 10043 350370
rect 9838 345491 10043 345692
rect 9838 345354 10038 345491
rect 9969 338749 10081 340759
rect 9969 338647 9974 338749
rect 10076 338647 10081 338749
rect 9969 338642 10081 338647
rect 9974 338638 10076 338642
rect 15780 305840 15880 509937
rect 18316 508772 18325 508972
rect 18525 508772 18534 508972
rect 9935 305740 15880 305840
rect 9935 302703 10035 305740
rect 9873 302332 10073 302703
rect 9953 295527 10065 297812
rect 9953 295425 9958 295527
rect 10060 295425 10065 295527
rect 9953 295420 10065 295425
rect 9958 295416 10060 295420
rect 18325 288719 18525 508772
rect 20797 488145 20806 488345
rect 21006 488145 21015 488345
rect 9889 288519 18525 288719
rect 9889 259222 10089 288519
rect 9956 252505 10068 254785
rect 9952 252403 9961 252505
rect 10063 252403 10072 252505
rect 9956 252398 10068 252403
rect 20806 241646 21006 488145
rect 9908 241446 21006 241646
rect 2293 214412 5870 214422
rect 2293 210749 5870 210759
rect 9908 131511 10108 241446
rect 9938 124883 10050 126976
rect 9938 124781 9943 124883
rect 10045 124781 10050 124883
rect 9938 124776 10050 124781
rect 9943 124772 10045 124776
rect 23823 116993 24023 543501
rect 430390 540770 430450 540779
rect 430390 540701 430450 540710
rect 26933 540436 26942 540636
rect 27142 540436 27151 540636
rect 9907 116793 24023 116993
rect 9907 88320 10107 116793
rect 9956 81661 10068 83810
rect 9952 81559 9961 81661
rect 10063 81559 10072 81661
rect 9956 81554 10068 81559
rect 26942 72999 27142 540436
rect 430397 538699 430443 540701
rect 430634 540423 430680 544234
rect 430934 540609 430980 544989
rect 437448 540735 437454 540830
rect 437549 540735 437555 540830
rect 430925 540557 430931 540609
rect 430983 540557 430989 540609
rect 430625 540371 430631 540423
rect 430683 540371 430689 540423
rect 437010 539801 437016 539888
rect 437103 539801 437109 539888
rect 433170 539495 433176 539600
rect 433281 539495 433287 539600
rect 430381 538639 430390 538699
rect 430450 538639 430459 538699
rect 30007 506074 30016 506274
rect 30216 506074 30225 506274
rect 9895 72799 27142 72999
rect 9895 44896 10095 72799
rect 9934 38439 10046 40414
rect 9934 38337 9939 38439
rect 10041 38337 10046 38439
rect 9934 38332 10046 38337
rect 9939 38328 10041 38332
rect 30016 34966 30216 506074
rect 433176 488245 433281 539495
rect 433167 488140 433176 488245
rect 433281 488140 433290 488245
rect 437016 480678 437103 539801
rect 437454 481879 437548 540735
rect 438114 534851 438204 546902
rect 438596 544475 438684 544481
rect 447254 544409 447300 555319
rect 447422 544531 447468 555576
rect 447413 544479 447419 544531
rect 447471 544479 447477 544531
rect 438596 535404 438684 544387
rect 447251 544403 447303 544409
rect 447251 544345 447303 544351
rect 439079 541783 439085 541900
rect 439202 541783 439208 541900
rect 439085 535886 439202 541783
rect 439817 541357 439823 541438
rect 439904 541357 439910 541438
rect 439542 541127 439548 541223
rect 439644 541127 439650 541223
rect 439548 536533 439644 541127
rect 439823 536999 439904 541357
rect 440096 541065 440181 541071
rect 440096 537343 440181 540980
rect 447176 539576 447236 539582
rect 440537 538965 440543 539052
rect 440630 538965 440636 539052
rect 440078 537268 440087 537343
rect 440189 537268 440198 537343
rect 440096 537263 440181 537268
rect 439814 536918 439823 536999
rect 439904 536918 439913 536999
rect 439539 536437 439548 536533
rect 439644 536437 439653 536533
rect 439085 535760 439202 535769
rect 438587 535316 438596 535404
rect 438684 535316 438693 535404
rect 438105 534761 438114 534851
rect 438204 534761 438213 534851
rect 437445 481785 437454 481879
rect 437548 481785 437557 481879
rect 437007 480591 437016 480678
rect 437103 480591 437112 480678
rect 440543 479746 440630 538965
rect 447176 538697 447236 539516
rect 447169 538641 447178 538697
rect 447234 538641 447243 538697
rect 447176 538639 447236 538641
rect 457047 529317 457147 555913
rect 458097 529803 459001 556700
rect 458097 529573 458416 529803
rect 458646 529573 459001 529803
rect 458097 529284 459001 529573
rect 457047 529208 457147 529217
rect 463400 528357 463800 556356
rect 482919 547053 482965 555882
rect 483341 555237 483387 555878
rect 483341 555191 483544 555237
rect 483498 547736 483544 555191
rect 483495 547730 483547 547736
rect 483495 547672 483547 547678
rect 482916 547047 482968 547053
rect 482916 546989 482968 546995
rect 576957 537348 577069 585931
rect 576948 537236 576957 537348
rect 577069 537236 577078 537348
rect 576981 536994 577062 536999
rect 576977 536923 576986 536994
rect 577057 536923 577066 536994
rect 575729 536528 575825 536533
rect 575725 536442 575734 536528
rect 575820 536442 575829 536528
rect 574240 535881 574357 535886
rect 574236 535774 574245 535881
rect 574352 535774 574361 535881
rect 572959 535404 573037 535408
rect 572954 535399 573042 535404
rect 572954 535321 572959 535399
rect 573037 535321 573042 535399
rect 571943 534846 572033 534851
rect 571939 534766 571948 534846
rect 572028 534766 572037 534846
rect 463391 527957 463400 528357
rect 463800 527957 463809 528357
rect 567420 489123 567429 489235
rect 567541 489123 567550 489235
rect 440534 479659 440543 479746
rect 440630 479659 440639 479746
rect 567429 269337 567541 489123
rect 571943 316101 572033 534766
rect 572954 361339 573042 535321
rect 574240 407799 574357 535774
rect 575729 452183 575825 536442
rect 576981 496608 577062 536923
rect 576972 496527 576981 496608
rect 577062 496527 577071 496608
rect 575720 452087 575729 452183
rect 575825 452087 575834 452183
rect 574231 407682 574240 407799
rect 574357 407682 574366 407799
rect 572945 361251 572954 361339
rect 573042 361251 573051 361339
rect 571934 316011 571943 316101
rect 572033 316011 572042 316101
rect 567425 269235 567434 269337
rect 567536 269235 567545 269337
rect 567429 269230 567541 269235
rect 253542 235028 253598 235047
rect 253542 234972 253861 235028
rect 253542 234936 253598 234972
rect 252906 233405 252978 233414
rect 203019 233398 203080 233401
rect 203012 233342 203021 233398
rect 203077 233342 203086 233398
rect 203019 124478 203080 233342
rect 252978 233383 253296 233405
rect 252978 233355 253584 233383
rect 252978 233333 253296 233355
rect 252906 233324 252978 233333
rect 253805 232982 253861 234972
rect 316562 234840 317290 234896
rect 317234 233706 317290 234840
rect 380379 234115 381167 234132
rect 379596 234087 381167 234115
rect 380379 234070 381167 234087
rect 381229 234070 381238 234132
rect 415039 234129 415101 234132
rect 415033 234073 415042 234129
rect 415098 234073 415107 234129
rect 318256 233706 318265 233708
rect 317234 233650 318265 233706
rect 317234 233603 317290 233650
rect 318256 233648 318265 233650
rect 318325 233648 318334 233708
rect 204294 213184 204404 213188
rect 204289 213179 204409 213184
rect 204289 213069 204294 213179
rect 204404 213069 204409 213179
rect 204289 212732 204409 213069
rect 9856 34766 30216 34966
rect 197880 124417 203080 124478
rect 9856 23515 10056 34766
rect 9944 17017 10055 19039
rect 9940 16916 9949 17017
rect 10050 16916 10059 17017
rect 9944 16911 10055 16916
rect 197880 8377 197941 124417
rect 204322 122655 204376 212732
rect 411942 188019 412062 188024
rect 411938 187909 411947 188019
rect 412057 187909 412066 188019
rect 411942 187477 412062 187909
rect 411965 186732 412040 187477
rect 411965 186657 413237 186732
rect 192883 8316 197941 8377
rect 201147 122601 204376 122655
rect 192883 3036 192944 8316
rect 201147 4489 201201 122601
rect 203449 120019 203569 120024
rect 203445 119909 203454 120019
rect 203564 119909 203573 120019
rect 203449 119663 203569 119909
rect 198164 4435 201201 4489
rect 192883 2975 194463 3036
rect 194402 480 194463 2975
rect 198164 1534 198218 4435
rect 203484 2067 203535 119663
rect 411762 94615 411882 94620
rect 411758 94505 411767 94615
rect 411877 94505 411886 94615
rect 411762 94193 411882 94505
rect 268276 26946 268586 26974
rect 205242 2082 205298 26170
rect 203484 2016 203919 2067
rect 205242 2026 208633 2082
rect 197953 1480 198218 1534
rect 197953 480 198007 1480
rect 203868 480 203919 2016
rect 208577 480 208633 2026
rect 268558 1372 268586 26946
rect 331296 26926 331547 26954
rect 394316 26932 394617 26960
rect 268558 1344 268909 1372
rect 268881 480 268909 1344
rect 331519 480 331547 26926
rect 394589 1932 394617 26932
rect 394589 1904 395371 1932
rect 395343 1122 395371 1904
rect 411779 1433 411866 94193
rect 413162 1845 413237 186657
rect 415039 2374 415101 234073
rect 415825 233706 415885 233708
rect 415818 233650 415827 233706
rect 415883 233650 415892 233706
rect 415825 10536 415885 233650
rect 415816 10476 415825 10536
rect 415885 10476 415894 10536
rect 579737 10534 579797 10536
rect 579730 10478 579739 10534
rect 579795 10478 579804 10534
rect 415039 2312 421398 2374
rect 413162 1770 416675 1845
rect 411779 1346 413141 1433
rect 395343 1094 396565 1122
rect 395343 1088 395371 1094
rect 396537 480 396565 1094
rect 413054 480 413141 1346
rect 416600 480 416675 1770
rect 421336 480 421398 2312
rect 579737 480 579797 10478
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 170994 700500 172994 701000
rect 222694 700500 224694 701000
rect 324394 700500 326394 701000
rect 576962 585931 577064 586033
rect 446236 548061 446814 549540
rect 430909 545043 430987 545121
rect 430628 544276 430684 544332
rect 23823 543501 24023 543701
rect 5911 537274 8454 541333
rect 8454 537274 9970 541333
rect 11305 523081 11555 523331
rect 6825 509177 6919 509271
rect 6830 481790 6914 481874
rect 5296 480596 5373 480673
rect 3076 479664 3153 479741
rect 5291 465976 5378 466063
rect 3071 422737 3158 422824
rect 15785 509937 15875 510027
rect 13411 507720 13601 507910
rect 11300 381827 11560 382087
rect 9974 338647 10076 338749
rect 18325 508772 18525 508972
rect 9958 295425 10060 295527
rect 20806 488145 21006 488345
rect 9961 252403 10063 252505
rect 2293 210759 5870 214412
rect 9943 124781 10045 124883
rect 430390 540710 430450 540770
rect 26942 540436 27142 540636
rect 9961 81559 10063 81661
rect 430390 538639 430450 538699
rect 30016 506074 30216 506274
rect 9939 38337 10041 38439
rect 433176 488140 433281 488245
rect 441536 539379 441976 540459
rect 440087 537268 440189 537343
rect 439823 536918 439904 536999
rect 439548 536437 439644 536533
rect 439085 535769 439202 535886
rect 438596 535316 438684 535404
rect 438114 534761 438204 534851
rect 437454 481785 437548 481879
rect 437016 480591 437103 480678
rect 447178 538641 447234 538697
rect 457047 529217 457147 529317
rect 458416 529573 458646 529803
rect 576957 537236 577069 537348
rect 576986 536923 577057 536994
rect 575734 536442 575820 536528
rect 574245 535774 574352 535881
rect 572959 535321 573037 535399
rect 571948 534766 572028 534846
rect 463400 527957 463800 528357
rect 567429 489123 567541 489235
rect 440543 479659 440630 479746
rect 576981 496527 577062 496608
rect 575729 452087 575825 452183
rect 574240 407682 574357 407799
rect 572954 361251 573042 361339
rect 571943 316011 572033 316101
rect 567434 269235 567536 269337
rect 203021 233342 203077 233398
rect 252906 233333 252978 233405
rect 381167 234070 381229 234132
rect 415042 234073 415098 234129
rect 318265 233648 318325 233708
rect 204294 213069 204404 213179
rect 9949 16916 10050 17017
rect 411947 187909 412057 188019
rect 203454 119909 203564 120019
rect 411767 94505 411877 94615
rect 415827 233650 415883 233706
rect 415825 10476 415885 10536
rect 579739 10478 579795 10534
<< metal3 >>
rect 16194 702200 21194 704800
rect 16194 701400 16294 702200
rect 21094 701400 21194 702200
rect 16194 701300 21194 701400
rect 16194 701000 21194 701100
rect 16194 700514 16294 701000
rect 3519 700200 16294 700514
rect 21094 700514 21194 701000
rect 68194 702200 73194 704800
rect 68194 701400 68294 702200
rect 73094 701400 73194 702200
rect 68194 701300 73194 701400
rect 68194 701000 73194 701100
rect 68194 700514 68294 701000
rect 21094 700200 68294 700514
rect 73094 700514 73194 701000
rect 120194 702200 125194 704800
rect 120194 701400 120294 702200
rect 125094 701400 125194 702200
rect 120194 701300 125194 701400
rect 120194 701000 125194 701100
rect 120194 700514 120294 701000
rect 73094 700200 120294 700514
rect 125094 700514 125194 701000
rect 165594 702200 170594 704800
rect 165594 701400 165694 702200
rect 170494 701400 170594 702200
rect 165594 701300 170594 701400
rect 165594 701000 170594 701100
rect 125094 700200 157105 700514
rect 3519 685242 157105 700200
rect -800 685142 2700 685242
rect -800 680342 1800 685142
rect 2600 680342 2700 685142
rect -800 680242 2700 680342
rect 2900 685142 157105 685242
rect 2900 680342 3000 685142
rect 3800 680342 157105 685142
rect 2900 680242 157105 680342
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect 3519 589976 157105 680242
rect 165594 700200 165694 701000
rect 170494 700200 170594 701000
rect 170894 701300 173094 704800
rect 170894 701000 173094 701100
rect 170894 700500 170994 701000
rect 172994 700500 173094 701000
rect 170894 700400 173094 700500
rect 173394 701300 175594 704800
rect 165594 700100 170594 700200
rect 173394 700100 175594 701100
rect 175894 702200 180894 704800
rect 175894 701400 175994 702200
rect 180794 701400 180894 702200
rect 175894 701300 180894 701400
rect 175894 701000 180894 701100
rect 175894 700200 175994 701000
rect 180794 700200 180894 701000
rect 175894 700100 180894 700200
rect 217294 702200 222294 704800
rect 217294 701400 217394 702200
rect 222194 701400 222294 702200
rect 217294 701300 222294 701400
rect 217294 701000 222294 701100
rect 217294 700200 217394 701000
rect 222194 700200 222294 701000
rect 222594 701300 224794 704800
rect 222594 701000 224794 701100
rect 222594 700500 222694 701000
rect 224694 700500 224794 701000
rect 222594 700400 224794 700500
rect 225094 701300 227294 704800
rect 217294 700100 222294 700200
rect 225094 700100 227294 701100
rect 227594 702200 232594 704800
rect 227594 701400 227694 702200
rect 232494 701400 232594 702200
rect 227594 701300 232594 701400
rect 227594 701000 232594 701100
rect 227594 700200 227694 701000
rect 232494 700200 232594 701000
rect 227594 700100 232594 700200
rect 318994 702200 323994 704800
rect 318994 701400 319094 702200
rect 323894 701400 323994 702200
rect 318994 701300 323994 701400
rect 318994 701000 323994 701100
rect 318994 700200 319094 701000
rect 323894 700200 323994 701000
rect 324294 701300 326494 704800
rect 324294 701000 326494 701100
rect 324294 700500 324394 701000
rect 326394 700500 326494 701000
rect 324294 700400 326494 700500
rect 326794 701300 328994 704800
rect 318994 700100 323994 700200
rect 326794 700100 328994 701100
rect 329294 702200 334294 704800
rect 329294 701400 329394 702200
rect 334194 701400 334294 702200
rect 329294 701300 334294 701400
rect 329294 701000 334294 701100
rect 329294 700200 329394 701000
rect 334194 700200 334294 701000
rect 329294 700100 334294 700200
rect 413394 702200 418394 704800
rect 413394 701400 413494 702200
rect 418294 701400 418394 702200
rect 413394 701300 418394 701400
rect 413394 701000 418394 701100
rect 413394 700200 413494 701000
rect 418294 700200 418394 701000
rect 413394 700100 418394 700200
rect 465394 702200 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 465394 701400 465494 702200
rect 470294 701400 470394 702200
rect 465394 701300 470394 701400
rect 465394 701000 470394 701100
rect 465394 700200 465494 701000
rect 470294 700200 470394 701000
rect 465394 700100 470394 700200
rect 566594 702200 571594 704800
rect 566594 701400 566694 702200
rect 571494 701400 571594 702200
rect 566594 701300 571594 701400
rect 566594 701000 571594 701100
rect 566594 700200 566694 701000
rect 571494 700200 571594 701000
rect 566594 700100 571594 700200
rect 165594 686800 384400 700100
rect 388400 686800 571594 700100
rect 165594 596000 344400 686800
rect 582300 682982 584800 682984
rect 527700 682882 581100 682982
rect 527700 678082 580200 682882
rect 581000 678082 581100 682882
rect 527700 677982 581100 678082
rect 581300 682882 584800 682982
rect 581300 678082 581400 682882
rect 582200 678082 584800 682882
rect 581300 677984 584800 678082
rect 581300 677982 582300 677984
rect 527700 661200 580100 677982
rect 573611 643784 584800 644584
rect 572401 630564 572411 643784
rect 580740 639784 584800 643784
rect 580740 634584 582340 639784
rect 580740 630564 584800 634584
rect 573611 629784 584800 630564
rect 573611 629764 582340 629784
rect 3470 568431 378401 589976
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 576957 586033 584800 586038
rect 576957 585931 576962 586033
rect 577064 585931 584800 586033
rect 576957 585926 584800 585931
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 564238 1660 564242
rect -800 559442 6204 564238
rect 1466 558151 6204 559442
rect 1464 554242 6206 558151
rect 16311 556000 378401 568431
rect -800 549785 6206 554242
rect 582340 550562 584800 555362
rect -800 549442 14440 549785
rect 1464 544527 14440 549442
rect 446176 549540 446874 549600
rect 446176 548061 446236 549540
rect 446814 548061 446874 549540
rect 446176 548001 446874 548061
rect 1464 540877 4962 544527
rect 4961 535050 4962 540877
rect 14439 535050 14440 544527
rect 397112 546102 400812 546302
rect 23818 543701 24028 543706
rect 397112 543701 397312 546102
rect 23818 543501 23823 543701
rect 24023 543501 397312 543701
rect 398857 545534 400709 545734
rect 23818 543496 24028 543501
rect 398857 542570 399057 545534
rect 430537 545121 430992 545126
rect 430537 545043 430909 545121
rect 430987 545043 430992 545121
rect 430537 545038 430992 545043
rect 430623 544334 430689 544337
rect 430532 544332 430689 544334
rect 430532 544276 430628 544332
rect 430684 544276 430689 544332
rect 430532 544274 430689 544276
rect 430623 544271 430689 544274
rect 395507 542370 399057 542570
rect 26937 540636 27147 540641
rect 395507 540636 395707 542370
rect 430385 540770 430455 540775
rect 430328 540710 430390 540770
rect 430450 540710 430455 540770
rect 430385 540705 430455 540710
rect 26937 540436 26942 540636
rect 27142 540436 395707 540636
rect 582340 540562 584800 545362
rect 441476 540459 442036 540519
rect 26937 540431 27147 540436
rect 441476 539379 441536 540459
rect 441976 539379 442036 540459
rect 441476 539319 442036 539379
rect 430385 538699 430455 538704
rect 447173 538699 447239 538702
rect 430385 538639 430390 538699
rect 430450 538697 447239 538699
rect 430450 538641 447178 538697
rect 447234 538641 447239 538697
rect 430450 538639 447239 538641
rect 430385 538634 430455 538639
rect 447173 538636 447239 538639
rect 576952 537348 577074 537353
rect 440082 537343 576957 537348
rect 440082 537268 440087 537343
rect 440189 537268 576957 537343
rect 440082 537236 576957 537268
rect 577069 537236 577074 537348
rect 576952 537231 577074 537236
rect 439818 536999 439909 537004
rect 439818 536918 439823 536999
rect 439904 536994 577062 536999
rect 439904 536923 576986 536994
rect 577057 536923 577062 536994
rect 439904 536918 577062 536923
rect 439818 536913 439909 536918
rect 439543 536533 439649 536538
rect 439543 536437 439548 536533
rect 439644 536528 575825 536533
rect 439644 536442 575734 536528
rect 575820 536442 575825 536528
rect 439644 536437 575825 536442
rect 439543 536432 439649 536437
rect 439080 535886 439207 535891
rect 439080 535769 439085 535886
rect 439202 535881 574357 535886
rect 439202 535774 574245 535881
rect 574352 535774 574357 535881
rect 439202 535769 574357 535774
rect 439080 535764 439207 535769
rect 438591 535404 438689 535409
rect 438591 535316 438596 535404
rect 438684 535399 573042 535404
rect 438684 535321 572959 535399
rect 573037 535321 573042 535399
rect 438684 535316 573042 535321
rect 438591 535311 438689 535316
rect 4961 535049 14440 535050
rect 4962 535044 14439 535049
rect 438109 534851 438209 534856
rect 438109 534761 438114 534851
rect 438204 534846 572033 534851
rect 438204 534766 571948 534846
rect 572028 534766 572033 534846
rect 438204 534761 572033 534766
rect 438109 534756 438209 534761
rect 430581 529803 458651 529808
rect 430581 529573 458416 529803
rect 458646 529573 458651 529803
rect 430581 529568 458651 529573
rect 430844 529317 431642 529370
rect 457042 529317 457152 529322
rect 430844 529270 457047 529317
rect 431542 529217 457047 529270
rect 457147 529217 457152 529317
rect 457042 529212 457152 529217
rect 430742 528936 431245 529036
rect 431145 528515 431245 528936
rect 431145 528415 462316 528515
rect 462216 528196 462316 528415
rect 463395 528357 463805 528362
rect 463395 528196 463400 528357
rect 462216 528096 463400 528196
rect 463395 527957 463400 528096
rect 463800 527957 463805 528357
rect 463395 527952 463805 527957
rect 11300 523331 401109 523336
rect 11300 523081 11305 523331
rect 11555 523081 401109 523331
rect 11300 523076 401109 523081
rect -800 511530 480 511642
rect -800 510348 480 510460
rect 15780 510027 400330 510032
rect 15780 509937 15785 510027
rect 15875 509937 400330 510027
rect 15780 509932 400330 509937
rect -800 509271 480 509278
rect 6820 509271 6924 509276
rect -800 509177 6825 509271
rect 6919 509177 6924 509271
rect -800 509166 480 509177
rect 6820 509172 6924 509177
rect 18320 508972 18530 508977
rect 18320 508772 18325 508972
rect 18525 508929 398631 508972
rect 18525 508829 399179 508929
rect 18525 508772 398631 508829
rect 18320 508767 18530 508772
rect 399079 508196 399179 508829
rect 400230 508441 400330 509932
rect 400230 508341 400746 508441
rect 399079 508096 400748 508196
rect -800 507984 480 508096
rect 13406 507910 400827 507915
rect 13406 507720 13411 507910
rect 13601 507720 400827 507910
rect 13406 507715 400827 507720
rect -800 506802 480 506914
rect 30011 506274 30221 506279
rect 30011 506074 30016 506274
rect 30216 506074 398321 506274
rect 30011 506069 30221 506074
rect -800 505620 480 505732
rect 398121 505520 398321 506074
rect 398121 505320 400866 505520
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 576976 496608 577067 496613
rect 583520 496608 584800 496616
rect 576976 496527 576981 496608
rect 577062 496527 584800 496608
rect 576976 496522 577067 496527
rect 583520 496504 584800 496527
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 567424 489235 567546 489240
rect 431956 489123 567429 489235
rect 567541 489123 567546 489235
rect 431956 488998 432068 489123
rect 567424 489118 567546 489123
rect 430675 488886 432068 488998
rect 20801 488345 21011 488350
rect 20801 488145 20806 488345
rect 21006 488145 406951 488345
rect 433171 488245 433286 488250
rect 20801 488140 21011 488145
rect 430394 488140 433176 488245
rect 433281 488140 433286 488245
rect 433171 488135 433286 488140
rect 437449 481879 437553 481884
rect 6825 481874 437454 481879
rect 6825 481790 6830 481874
rect 6914 481790 437454 481874
rect 6825 481785 437454 481790
rect 437548 481785 437553 481879
rect 437449 481780 437553 481785
rect 437011 480678 437108 480683
rect 5291 480673 437016 480678
rect 5291 480596 5296 480673
rect 5373 480596 437016 480673
rect 5291 480591 437016 480596
rect 437103 480591 437108 480678
rect 437011 480586 437108 480591
rect 440538 479746 440635 479751
rect 3071 479741 440543 479746
rect 3071 479664 3076 479741
rect 3153 479664 440543 479741
rect 3071 479659 440543 479664
rect 440630 479659 440635 479746
rect 440538 479654 440635 479659
rect -800 468308 480 468420
rect -800 467126 480 467238
rect 5286 466063 5383 466068
rect 272 466056 5291 466063
rect -800 465976 5291 466056
rect 5378 465976 5383 466063
rect -800 465944 480 465976
rect 5286 465971 5383 465976
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 575724 452183 575830 452188
rect 583520 452183 584800 452194
rect 575724 452087 575729 452183
rect 575825 452087 584800 452183
rect 575724 452082 575830 452087
rect 583520 452082 584800 452087
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422824 480 422834
rect 3066 422824 3163 422829
rect -800 422737 3071 422824
rect 3158 422737 3163 422824
rect -800 422722 480 422737
rect 3066 422732 3163 422737
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 574235 407799 574362 407804
rect 574235 407682 574240 407799
rect 574357 407772 583772 407799
rect 574357 407682 584800 407772
rect 574235 407677 574362 407682
rect 583520 407660 584800 407682
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 11295 382087 11565 382092
rect 11038 382062 11300 382087
rect 875 381976 11300 382062
rect -800 381864 11300 381976
rect 875 381827 11300 381864
rect 11560 381827 11565 382087
rect 875 381822 11565 381827
rect 875 381802 11499 381822
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 572949 361339 573047 361344
rect 583520 361339 584800 361350
rect 572949 361251 572954 361339
rect 573042 361251 584800 361339
rect 572949 361246 573047 361251
rect 583520 361238 584800 361251
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338749 10081 338754
rect -800 338647 9974 338749
rect 10076 338647 10081 338749
rect -800 338642 10081 338647
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 571938 316101 572038 316106
rect 583520 316101 584800 316128
rect 571938 316011 571943 316101
rect 572033 316016 584800 316101
rect 572033 316011 583667 316016
rect 571938 316006 572038 316011
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295527 10065 295532
rect -800 295425 9958 295527
rect 10060 295425 10065 295527
rect -800 295420 10065 295425
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 567429 269337 584800 269342
rect 567429 269235 567434 269337
rect 567536 269235 584800 269337
rect 567429 269230 584800 269235
rect -800 252505 10068 252510
rect -800 252403 9961 252505
rect 10063 252403 10068 252505
rect -800 252398 10068 252403
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 381162 234132 381234 234137
rect 415037 234132 415103 234134
rect 381162 234070 381167 234132
rect 381229 234129 415103 234132
rect 381229 234073 415042 234129
rect 415098 234073 415103 234129
rect 381229 234070 415103 234073
rect 381162 234065 381234 234070
rect 415037 234068 415103 234070
rect 318260 233708 318330 233713
rect 415822 233708 415888 233711
rect 318260 233648 318265 233708
rect 318325 233706 415888 233708
rect 318325 233650 415827 233706
rect 415883 233650 415888 233706
rect 318325 233648 415888 233650
rect 318260 233643 318330 233648
rect 415822 233645 415888 233648
rect 252901 233405 252983 233410
rect 203016 233400 203082 233403
rect 252494 233400 252906 233405
rect 203016 233398 252906 233400
rect 203016 233342 203021 233398
rect 203077 233342 252906 233398
rect 203016 233339 252906 233342
rect 203016 233337 203082 233339
rect 252494 233333 252906 233339
rect 252978 233333 252983 233405
rect 252901 233328 252983 233333
rect 582340 225230 584800 230030
rect 1229 219889 17420 220141
rect 1229 219688 4477 219889
rect -800 214888 4477 219688
rect 1229 214412 4477 214888
rect 1229 210759 2293 214412
rect 1229 210412 4477 210759
rect 13954 210412 17420 219889
rect 204289 213179 204884 213184
rect 204289 213069 204294 213179
rect 204404 213069 204884 213179
rect 204289 213064 204884 213069
rect 1229 209688 17420 210412
rect -800 204888 17420 209688
rect 1229 204791 17420 204888
rect 572045 195230 584800 196230
rect 411436 188019 412062 188024
rect 411436 187909 411947 188019
rect 412057 187909 412062 188019
rect 411436 187904 412062 187909
rect 572045 182430 573045 195230
rect 580340 191430 584800 195230
rect 580340 186230 582340 191430
rect 580340 182430 584800 186230
rect 572045 181430 584800 182430
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124883 10050 124888
rect -800 124781 9943 124883
rect 10045 124781 10050 124883
rect -800 124776 10050 124781
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect 203858 120024 203976 120029
rect 203449 120023 203977 120024
rect 203449 120019 203858 120023
rect 203449 119909 203454 120019
rect 203564 119909 203858 120019
rect 203449 119905 203858 119909
rect 203976 119905 203977 120023
rect 203449 119904 203977 119905
rect 204294 119904 204300 120024
rect 204420 119904 204884 120024
rect 203858 119899 203976 119904
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 411436 94744 411882 94864
rect 411762 94615 411882 94744
rect 411762 94505 411767 94615
rect 411877 94505 411882 94615
rect 411762 94500 411882 94505
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81661 10068 81666
rect -800 81559 9961 81661
rect 10063 81559 10068 81661
rect -800 81554 10068 81559
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38439 10046 38444
rect -800 38337 9939 38439
rect 10041 38337 10046 38439
rect -800 38332 10046 38337
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 17017 10055 17022
rect -800 16916 9949 17017
rect 10050 16916 10055 17017
rect -800 16911 10055 16916
rect -800 16910 480 16911
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect 415820 10536 415890 10541
rect 579734 10536 579800 10539
rect 415820 10476 415825 10536
rect 415885 10534 579800 10536
rect 415885 10478 579739 10534
rect 579795 10478 579800 10534
rect 415885 10476 579800 10478
rect 415820 10471 415890 10476
rect 579734 10473 579800 10476
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 16194 701100 21194 701300
rect 68194 701100 73194 701300
rect 120194 701100 125194 701300
rect 165594 701100 170594 701300
rect 2700 680242 2900 685242
rect 170894 701100 173094 701300
rect 173394 701100 175594 701300
rect 175894 701100 180894 701300
rect 217294 701100 222294 701300
rect 222594 701100 224794 701300
rect 225094 701100 227294 701300
rect 227594 701100 232594 701300
rect 318994 701100 323994 701300
rect 324294 701100 326494 701300
rect 326794 701100 328994 701300
rect 329294 701100 334294 701300
rect 413394 701100 418394 701300
rect 465394 701100 470394 701300
rect 566594 701100 571594 701300
rect 581100 677982 581300 682982
<< via3 >>
rect 16294 701400 21094 702200
rect 16294 700200 21094 701000
rect 68294 701400 73094 702200
rect 68294 700200 73094 701000
rect 120294 701400 125094 702200
rect 120294 700200 125094 701000
rect 165694 701400 170494 702200
rect 1800 680342 2600 685142
rect 3000 680342 3800 685142
rect 165694 700200 170494 701000
rect 175994 701400 180794 702200
rect 175994 700200 180794 701000
rect 217394 701400 222194 702200
rect 217394 700200 222194 701000
rect 227694 701400 232494 702200
rect 227694 700200 232494 701000
rect 319094 701400 323894 702200
rect 319094 700200 323894 701000
rect 329394 701400 334194 702200
rect 329394 700200 334194 701000
rect 413494 701400 418294 702200
rect 413494 700200 418294 701000
rect 465494 701400 470294 702200
rect 465494 700200 470294 701000
rect 566694 701400 571494 702200
rect 566694 700200 571494 701000
rect 580200 678082 581000 682882
rect 581400 678082 582200 682882
rect 572411 630564 580740 643784
rect 446236 548061 446814 549540
rect 4962 541333 14439 544527
rect 4962 537274 5911 541333
rect 5911 537274 9970 541333
rect 9970 537274 14439 541333
rect 4962 535050 14439 537274
rect 441536 539379 441976 540459
rect 4477 214412 13954 219889
rect 4477 210759 5870 214412
rect 5870 210759 13954 214412
rect 4477 210412 13954 210759
rect 573045 182430 580340 195230
rect 203858 119905 203976 120023
rect 204300 119904 204420 120024
<< metal4 >>
rect 16194 702200 21194 702300
rect 16194 701400 16294 702200
rect 21094 701400 21194 702200
rect 16194 701300 21194 701400
rect 16194 701000 21194 701100
rect 16194 700514 16294 701000
rect 3519 700200 16294 700514
rect 21094 700514 21194 701000
rect 68194 702200 73194 702300
rect 68194 701400 68294 702200
rect 73094 701400 73194 702200
rect 68194 701300 73194 701400
rect 68194 701000 73194 701100
rect 68194 700514 68294 701000
rect 21094 700200 68294 700514
rect 73094 700514 73194 701000
rect 120194 702200 125194 702300
rect 120194 701400 120294 702200
rect 125094 701400 125194 702200
rect 120194 701300 125194 701400
rect 120194 701000 125194 701100
rect 120194 700514 120294 701000
rect 73094 700200 120294 700514
rect 125094 700514 125194 701000
rect 165594 702200 170594 702300
rect 165594 701400 165694 702200
rect 170494 701400 170594 702200
rect 165594 701300 170594 701400
rect 165594 701000 170594 701100
rect 125094 700200 157105 700514
rect 3519 685242 157105 700200
rect 1700 685142 2700 685242
rect 1700 680342 1800 685142
rect 2600 680342 2700 685142
rect 1700 680242 2700 680342
rect 2900 685142 157105 685242
rect 2900 680342 3000 685142
rect 3800 680342 157105 685142
rect 2900 680242 157105 680342
rect 3519 589976 157105 680242
rect 165594 700200 165694 701000
rect 170494 700200 170594 701000
rect 165594 700100 170594 700200
rect 175894 702200 180894 702300
rect 175894 701400 175994 702200
rect 180794 701400 180894 702200
rect 175894 701300 180894 701400
rect 175894 701000 180894 701100
rect 175894 700200 175994 701000
rect 180794 700200 180894 701000
rect 175894 700100 180894 700200
rect 217294 702200 222294 702300
rect 217294 701400 217394 702200
rect 222194 701400 222294 702200
rect 217294 701300 222294 701400
rect 217294 701000 222294 701100
rect 217294 700200 217394 701000
rect 222194 700200 222294 701000
rect 217294 700100 222294 700200
rect 227594 702200 232594 702300
rect 227594 701400 227694 702200
rect 232494 701400 232594 702200
rect 227594 701300 232594 701400
rect 227594 701000 232594 701100
rect 227594 700200 227694 701000
rect 232494 700200 232594 701000
rect 227594 700100 232594 700200
rect 318994 702200 323994 702300
rect 318994 701400 319094 702200
rect 323894 701400 323994 702200
rect 318994 701300 323994 701400
rect 318994 701000 323994 701100
rect 318994 700200 319094 701000
rect 323894 700200 323994 701000
rect 318994 700100 323994 700200
rect 329294 702200 334294 702300
rect 329294 701400 329394 702200
rect 334194 701400 334294 702200
rect 329294 701300 334294 701400
rect 329294 701000 334294 701100
rect 329294 700200 329394 701000
rect 334194 700200 334294 701000
rect 329294 700100 334294 700200
rect 413394 702200 418394 702300
rect 413394 701400 413494 702200
rect 418294 701400 418394 702200
rect 413394 701300 418394 701400
rect 413394 701000 418394 701100
rect 413394 700200 413494 701000
rect 418294 700200 418394 701000
rect 413394 700100 418394 700200
rect 465394 702200 470394 702300
rect 465394 701400 465494 702200
rect 470294 701400 470394 702200
rect 465394 701300 470394 701400
rect 465394 701000 470394 701100
rect 465394 700200 465494 701000
rect 470294 700200 470394 701000
rect 465394 700100 470394 700200
rect 566594 702200 571594 702300
rect 566594 701400 566694 702200
rect 571494 701400 571594 702200
rect 566594 701300 571594 701400
rect 566594 701000 571594 701100
rect 566594 700200 566694 701000
rect 571494 700200 571594 701000
rect 566594 700100 571594 700200
rect 165594 686800 384400 700100
rect 388400 686800 571594 700100
rect 165594 596000 344400 686800
rect 527700 682882 581100 682982
rect 527700 678082 580200 682882
rect 581000 678082 581100 682882
rect 527700 677982 581100 678082
rect 581300 682882 582300 682982
rect 581300 678082 581400 682882
rect 582200 678082 582300 682882
rect 581300 677982 582300 678082
rect 527700 661200 580100 677982
rect 572410 643784 580741 643785
rect 572410 630564 572411 643784
rect 580740 630564 580741 643784
rect 572410 630563 580741 630564
rect 3519 568431 378401 589976
rect 16311 556000 378401 568431
rect 395963 549511 402412 549600
rect 395963 548137 396606 549511
rect 398010 548137 402412 549511
rect 395963 548000 402412 548137
rect 429320 549540 446953 549600
rect 429320 548061 446236 549540
rect 446814 548061 446953 549540
rect 429320 548000 446953 548061
rect 4961 544527 401120 544528
rect 4961 535050 4962 544527
rect 14439 535050 401120 544527
rect 428320 540460 442098 540600
rect 428320 539239 433094 540460
rect 434699 540459 442098 540460
rect 434699 539379 441536 540459
rect 441976 539379 442098 540459
rect 434699 539239 442098 539379
rect 428320 539000 442098 539239
rect 4961 535049 401120 535050
rect 396284 531522 402123 531600
rect 396284 530148 396619 531522
rect 398023 530148 402123 531522
rect 396284 530000 402123 530148
rect 428492 530000 434927 531600
rect 427886 522501 435183 522602
rect 427886 521280 433086 522501
rect 434691 521280 435183 522501
rect 427886 520999 435183 521280
rect 15731 513600 399172 517132
rect 15731 513512 402925 513600
rect 15731 512138 396627 513512
rect 398031 512138 402925 513512
rect 15731 512000 402925 512138
rect 15731 507653 399172 512000
rect 15731 219890 25210 507653
rect 428269 504417 435245 504600
rect 428269 503196 433127 504417
rect 434732 503196 435245 504417
rect 428269 503000 435245 503196
rect 397628 501200 409656 502000
rect 399806 493673 408961 493800
rect 399806 492308 399879 493673
rect 400615 492308 408961 493673
rect 399806 492200 408961 492308
rect 397684 484000 408654 484800
rect 208972 232424 209292 243254
rect 224332 232356 224652 234604
rect 239692 232424 240012 243106
rect 255052 232464 255372 234268
rect 270412 232424 270732 242828
rect 285772 232504 286092 234350
rect 301132 232422 301452 242868
rect 316492 232504 316812 235254
rect 331852 232424 332172 242656
rect 347212 232446 347532 234458
rect 362572 232424 362892 242812
rect 377932 232504 378252 234260
rect 393292 232424 393612 242754
rect 408652 232390 408972 234392
rect 4476 219889 25210 219890
rect 4476 210412 4477 219889
rect 13954 210412 25210 219889
rect 4476 210411 25210 210412
rect 573044 195230 580341 195231
rect 573044 182430 573045 195230
rect 580340 182430 580341 195230
rect 573044 182429 580341 182430
rect 204299 120024 204421 120025
rect 203857 120023 204300 120024
rect 203857 119905 203858 120023
rect 203976 119905 204300 120023
rect 203857 119904 204300 119905
rect 204420 119904 204421 120024
rect 204299 119903 204421 119904
<< rmetal4 >>
rect 16194 701100 21194 701300
rect 68194 701100 73194 701300
rect 120194 701100 125194 701300
rect 165594 701100 170594 701300
rect 2700 680242 2900 685242
rect 175894 701100 180894 701300
rect 217294 701100 222294 701300
rect 227594 701100 232594 701300
rect 318994 701100 323994 701300
rect 329294 701100 334294 701300
rect 413394 701100 418394 701300
rect 465394 701100 470394 701300
rect 566594 701100 571594 701300
rect 581100 677982 581300 682982
<< via4 >>
rect 16294 701400 21094 702200
rect 16294 700200 21094 701000
rect 68294 701400 73094 702200
rect 68294 700200 73094 701000
rect 120294 701400 125094 702200
rect 120294 700200 125094 701000
rect 165694 701400 170494 702200
rect 1800 680342 2600 685142
rect 3000 680342 3800 685142
rect 165694 700200 170494 701000
rect 175994 701400 180794 702200
rect 175994 700200 180794 701000
rect 217394 701400 222194 702200
rect 217394 700200 222194 701000
rect 227694 701400 232494 702200
rect 227694 700200 232494 701000
rect 319094 701400 323894 702200
rect 319094 700200 323894 701000
rect 329394 701400 334194 702200
rect 329394 700200 334194 701000
rect 413494 701400 418294 702200
rect 413494 700200 418294 701000
rect 465494 701400 470294 702200
rect 465494 700200 470294 701000
rect 566694 701400 571494 702200
rect 566694 700200 571494 701000
rect 580200 678082 581000 682882
rect 581400 678082 582200 682882
rect 572411 630564 580740 643784
rect 396606 548137 398010 549511
rect 433094 539239 434699 540460
rect 396619 530148 398023 531522
rect 433086 521280 434691 522501
rect 396627 512138 398031 513512
rect 433127 503196 434732 504417
rect 396828 501200 397628 502000
rect 399879 492308 400615 493673
rect 396884 484000 397684 484800
rect 208972 243254 209292 243574
rect 239692 243106 240012 243426
rect 224332 234604 224652 234924
rect 270412 242828 270732 243148
rect 255052 234268 255372 234588
rect 301132 242868 301452 243188
rect 285772 234350 286092 234670
rect 331852 242656 332172 242976
rect 316492 235254 316812 235574
rect 362572 242812 362892 243132
rect 347212 234458 347532 234778
rect 393292 242754 393612 243074
rect 377932 234260 378252 234580
rect 408652 234392 408972 234712
rect 573045 182430 580340 195230
<< metal5 >>
rect 16194 702200 21194 702300
rect 16194 701400 16294 702200
rect 21094 701400 21194 702200
rect 16194 701300 21194 701400
rect 16194 701000 21194 701100
rect 16194 700514 16294 701000
rect 3519 700200 16294 700514
rect 21094 700514 21194 701000
rect 68194 702200 73194 702300
rect 68194 701400 68294 702200
rect 73094 701400 73194 702200
rect 68194 701300 73194 701400
rect 68194 701000 73194 701100
rect 68194 700514 68294 701000
rect 21094 700200 68294 700514
rect 73094 700514 73194 701000
rect 120194 702200 125194 702300
rect 120194 701400 120294 702200
rect 125094 701400 125194 702200
rect 120194 701300 125194 701400
rect 120194 701000 125194 701100
rect 120194 700514 120294 701000
rect 73094 700200 120294 700514
rect 125094 700514 125194 701000
rect 165594 702200 170594 702300
rect 165594 701400 165694 702200
rect 170494 701400 170594 702200
rect 165594 701300 170594 701400
rect 165594 701000 170594 701100
rect 125094 700200 157105 700514
rect 3519 685242 157105 700200
rect 1700 685142 2700 685242
rect 1700 680342 1800 685142
rect 2600 680342 2700 685142
rect 1700 680242 2700 680342
rect 2900 685142 157105 685242
rect 2900 680342 3000 685142
rect 3800 680342 157105 685142
rect 2900 680242 157105 680342
rect 3519 589976 157105 680242
rect 165594 700200 165694 701000
rect 170494 700200 170594 701000
rect 165594 700100 170594 700200
rect 175894 702200 180894 702300
rect 175894 701400 175994 702200
rect 180794 701400 180894 702200
rect 175894 701300 180894 701400
rect 175894 701000 180894 701100
rect 175894 700200 175994 701000
rect 180794 700200 180894 701000
rect 175894 700100 180894 700200
rect 217294 702200 222294 702300
rect 217294 701400 217394 702200
rect 222194 701400 222294 702200
rect 217294 701300 222294 701400
rect 217294 701000 222294 701100
rect 217294 700200 217394 701000
rect 222194 700200 222294 701000
rect 217294 700100 222294 700200
rect 227594 702200 232594 702300
rect 227594 701400 227694 702200
rect 232494 701400 232594 702200
rect 227594 701300 232594 701400
rect 227594 701000 232594 701100
rect 227594 700200 227694 701000
rect 232494 700200 232594 701000
rect 227594 700100 232594 700200
rect 318994 702200 323994 702300
rect 318994 701400 319094 702200
rect 323894 701400 323994 702200
rect 318994 701300 323994 701400
rect 318994 701000 323994 701100
rect 318994 700200 319094 701000
rect 323894 700200 323994 701000
rect 318994 700100 323994 700200
rect 329294 702200 334294 702300
rect 329294 701400 329394 702200
rect 334194 701400 334294 702200
rect 329294 701300 334294 701400
rect 329294 701000 334294 701100
rect 329294 700200 329394 701000
rect 334194 700200 334294 701000
rect 329294 700100 334294 700200
rect 413394 702200 418394 702300
rect 413394 701400 413494 702200
rect 418294 701400 418394 702200
rect 413394 701300 418394 701400
rect 413394 701000 418394 701100
rect 413394 700200 413494 701000
rect 418294 700200 418394 701000
rect 413394 700100 418394 700200
rect 465394 702200 470394 702300
rect 465394 701400 465494 702200
rect 470294 701400 470394 702200
rect 465394 701300 470394 701400
rect 465394 701000 470394 701100
rect 465394 700200 465494 701000
rect 470294 700200 470394 701000
rect 465394 700100 470394 700200
rect 566594 702200 571594 702300
rect 566594 701400 566694 702200
rect 571494 701400 571594 702200
rect 566594 701300 571594 701400
rect 566594 701000 571594 701100
rect 566594 700200 566694 701000
rect 571494 700200 571594 701000
rect 566594 700100 571594 700200
rect 165594 686800 384400 700100
rect 388400 686800 571594 700100
rect 165594 596000 344400 686800
rect 527700 682882 581100 682982
rect 527700 678082 580200 682882
rect 581000 678082 581100 682882
rect 527700 677982 581100 678082
rect 581300 682882 582300 682982
rect 581300 678082 581400 682882
rect 582200 678082 582300 682882
rect 581300 677982 582300 678082
rect 527700 661200 580100 677982
rect 571611 643784 581540 644584
rect 571611 630564 572411 643784
rect 580740 630564 581540 643784
rect 571611 629764 581540 630564
rect 3152 568431 378376 589976
rect 16311 556000 378376 568431
rect 396506 549511 398144 549756
rect 396506 548137 396606 549511
rect 398010 548137 398144 549511
rect 396506 531522 398144 548137
rect 396506 530148 396619 531522
rect 398023 530148 398144 531522
rect 396506 513512 398144 530148
rect 396506 512138 396627 513512
rect 398031 512138 398144 513512
rect 396506 502000 398144 512138
rect 432950 540460 434923 549429
rect 432950 539239 433094 540460
rect 434699 539239 434923 540460
rect 432950 522501 434923 539239
rect 571621 529888 579950 629764
rect 432950 521280 433086 522501
rect 434691 521280 434923 522501
rect 396506 501200 396828 502000
rect 397628 501200 398144 502000
rect 396506 484800 398144 501200
rect 396506 484000 396884 484800
rect 397684 484000 398144 484800
rect 396506 483611 398144 484000
rect 399800 493673 400800 505541
rect 399800 492308 399879 493673
rect 400615 492308 400800 493673
rect 399800 483963 400800 492308
rect 430800 484042 431800 505658
rect 432950 504417 434923 521280
rect 432950 503196 433127 504417
rect 434732 503196 434923 504417
rect 432950 484147 434923 503196
rect 560020 521559 579950 529888
rect 560020 341085 568349 521559
rect 459092 332756 568349 341085
rect 459092 268551 467421 332756
rect 396651 260222 467421 268551
rect 396651 249346 404980 260222
rect 205238 243574 410704 249346
rect 205238 243254 208972 243574
rect 209292 243426 410704 243574
rect 209292 243254 239692 243426
rect 205238 243106 239692 243254
rect 240012 243188 410704 243426
rect 240012 243148 301132 243188
rect 240012 243106 270412 243148
rect 205238 242828 270412 243106
rect 270732 242868 301132 243148
rect 301452 243132 410704 243188
rect 301452 242976 362572 243132
rect 301452 242868 331852 242976
rect 270732 242828 331852 242868
rect 205238 242656 331852 242828
rect 332172 242812 362572 242976
rect 362892 243074 410704 243132
rect 362892 242812 393292 243074
rect 332172 242754 393292 242812
rect 393612 242754 410704 243074
rect 332172 242656 410704 242754
rect 205238 242536 410704 242656
rect 205174 235574 506191 240914
rect 205174 235254 316492 235574
rect 316812 235254 506191 235574
rect 205174 234924 506191 235254
rect 205174 234604 224332 234924
rect 224652 234778 506191 234924
rect 224652 234670 347212 234778
rect 224652 234604 285772 234670
rect 205174 234588 285772 234604
rect 205174 234268 255052 234588
rect 255372 234350 285772 234588
rect 286092 234458 347212 234670
rect 347532 234712 506191 234778
rect 347532 234580 408652 234712
rect 347532 234458 377932 234580
rect 286092 234350 377932 234458
rect 255372 234268 377932 234350
rect 205174 234260 377932 234268
rect 378252 234392 408652 234580
rect 408972 234392 410640 234712
rect 378252 234260 410640 234392
rect 205174 234104 410640 234260
rect 499989 195176 506191 234712
rect 559584 195230 581340 196230
rect 559584 195176 573045 195230
rect 499989 188974 573045 195176
rect 559584 182430 573045 188974
rect 580340 182430 581340 195230
rect 559584 181435 581340 182430
rect 572045 181430 581340 181435
<< rm5 >>
rect 16194 701100 21194 701300
rect 68194 701100 73194 701300
rect 120194 701100 125194 701300
rect 165594 701100 170594 701300
rect 2700 680242 2900 685242
rect 175894 701100 180894 701300
rect 217294 701100 222294 701300
rect 227594 701100 232594 701300
rect 318994 701100 323994 701300
rect 329294 701100 334294 701300
rect 413394 701100 418394 701300
rect 465394 701100 470394 701300
rect 566594 701100 571594 701300
rect 581100 677982 581300 682982
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use snproc  snproc_0
timestamp 1624430562
transform 1 0 204764 0 1 26056
box 0 0 206792 208936
use esd_cell  esd_cell_0
timestamp 1624430562
transform 0 -1 10000 1 0 21200
box -2400 -3178 2400 3178
use esd_cell  esd_cell_1
timestamp 1624430562
transform 0 -1 10000 1 0 42600
box -2400 -3178 2400 3178
use esd_cell  esd_cell_2
timestamp 1624430562
transform 0 -1 10000 1 0 86000
box -2400 -3178 2400 3178
use esd_cell  esd_cell_3
timestamp 1624430562
transform 0 -1 10000 1 0 129200
box -2400 -3178 2400 3178
use esd_cell  esd_cell_6
timestamp 1624430562
transform 0 -1 10000 1 0 343000
box -2400 -3178 2400 3178
use esd_cell  esd_cell_4
timestamp 1624430562
transform 0 -1 10000 1 0 300000
box -2400 -3178 2400 3178
use esd_cell  esd_cell_5
timestamp 1624430562
transform 0 -1 10000 1 0 257000
box -2400 -3178 2400 3178
use oscillator  oscillator_0
timestamp 1624430562
transform 1 0 418800 0 1 493000
box -12000 -9000 12000 9000
use power_stage  power_stage_0
timestamp 1624430562
transform 1 0 463600 0 1 620000
box -119200 -64204 96100 66802
use analog_subsystem  analog_subsystem_0
timestamp 1624430562
transform 1 0 418800 0 1 530800
box -19000 -27800 13000 18800
use switch_control  switch_control_0
timestamp 1624430562
transform 1 0 441400 0 1 538400
box -66 771 5538 8997
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal2 205242 26022 205298 26025 1 FreeSans 800 0 0 0 msg_from_snproc_available
flabel metal3 204690 119904 204695 120024 1 FreeSans 800 0 0 0 control_mode_data_in
flabel metal3 204695 213064 204706 213184 1 FreeSans 800 0 0 0 debug_bit_bottom_of_r1
flabel metal2 253805 232982 253861 232994 1 FreeSans 400 0 0 0 control_mode_data_out
flabel metal2 317234 233603 317290 233617 1 FreeSans 800 0 0 0 clock
flabel metal2 379842 234087 379853 234115 1 FreeSans 800 0 0 0 error_occured
flabel metal3 411610 187904 411654 188024 1 FreeSans 800 0 0 0 control_mode_execute
flabel metal3 411663 94744 411678 94864 1 FreeSans 800 0 0 0 assert_control_mode
flabel metal2 394589 26074 394617 26086 1 FreeSans 800 0 0 0 msg_to_snproc_full
flabel metal2 331519 26594 331547 26613 1 FreeSans 800 0 0 0 control_mode_clock
flabel metal2 268558 26287 268586 26315 1 FreeSans 800 0 0 0 debug_bit_bottom_of_ip
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
